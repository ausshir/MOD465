
//RX Filter 18'sd Multiplier Coefficients (headroom)
assign coef[  0] = -18'sd    195;
assign coef[  1] = -18'sd    201;
assign coef[  2] = -18'sd     49;
assign coef[  3] =  18'sd    155;
assign coef[  4] =  18'sd    261;
assign coef[  5] =  18'sd    175;
assign coef[  6] = -18'sd     54;
assign coef[  7] = -18'sd    267;
assign coef[  8] = -18'sd    302;
assign coef[  9] = -18'sd    115;
assign coef[ 10] =  18'sd    176;
assign coef[ 11] =  18'sd    366;
assign coef[ 12] =  18'sd    306;
assign coef[ 13] =  18'sd     19;
assign coef[ 14] = -18'sd    305;
assign coef[ 15] = -18'sd    434;
assign coef[ 16] = -18'sd    262;
assign coef[ 17] =  18'sd    108;
assign coef[ 18] =  18'sd    421;
assign coef[ 19] =  18'sd    450;
assign coef[ 20] =  18'sd    159;
assign coef[ 21] = -18'sd    256;
assign coef[ 22] = -18'sd    500;
assign coef[ 23] = -18'sd    389;
assign coef[ 24] =  18'sd      9;
assign coef[ 25] =  18'sd    409;
assign coef[ 26] =  18'sd    512;
assign coef[ 27] =  18'sd    228;
assign coef[ 28] = -18'sd    245;
assign coef[ 29] = -18'sd    546;
assign coef[ 30] = -18'sd    425;
assign coef[ 31] =  18'sd     57;
assign coef[ 32] =  18'sd    545;
assign coef[ 33] =  18'sd    637;
assign coef[ 34] =  18'sd    201;
assign coef[ 35] = -18'sd    488;
assign coef[ 36] = -18'sd    902;
assign coef[ 37] = -18'sd    648;
assign coef[ 38] =  18'sd    203;
assign coef[ 39] =  18'sd   1088;
assign coef[ 40] =  18'sd   1304;
assign coef[ 41] =  18'sd    534;
assign coef[ 42] = -18'sd    838;
assign coef[ 43] = -18'sd   1885;
assign coef[ 44] = -18'sd   1734;
assign coef[ 45] = -18'sd    239;
assign coef[ 46] =  18'sd   1771;
assign coef[ 47] =  18'sd   2915;
assign coef[ 48] =  18'sd   2170;
assign coef[ 49] = -18'sd    316;
assign coef[ 50] = -18'sd   3103;
assign coef[ 51] = -18'sd   4246;
assign coef[ 52] = -18'sd   2592;
assign coef[ 53] =  18'sd   1253;
assign coef[ 54] =  18'sd   5011;
assign coef[ 55] =  18'sd   6010;
assign coef[ 56] =  18'sd   2976;
assign coef[ 57] = -18'sd   2808;
assign coef[ 58] = -18'sd   7876;
assign coef[ 59] = -18'sd   8526;
assign coef[ 60] = -18'sd   3301;
assign coef[ 61] =  18'sd   5533;
assign coef[ 62] =  18'sd  12690;
assign coef[ 63] =  18'sd  12713;
assign coef[ 64] =  18'sd   3547;
assign coef[ 65] = -18'sd  11229;
assign coef[ 66] = -18'sd  23132;
assign coef[ 67] = -18'sd  22523;
assign coef[ 68] = -18'sd   3702;
assign coef[ 69] =  18'sd  31309;
assign coef[ 70] =  18'sd  72493;
assign coef[ 71] =  18'sd 105590;
assign coef[ 72] =  18'sd 118244;
