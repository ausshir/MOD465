
//RX Filter 18'sd Multiplier Coefficients (headroom)
assign coef[  0] = -18'sd     42;
assign coef[  1] =  18'sd     20;
assign coef[  2] =  18'sd     71;
assign coef[  3] =  18'sd     73;
assign coef[  4] =  18'sd     22;
assign coef[  5] = -18'sd     48;
assign coef[  6] = -18'sd     87;
assign coef[  7] = -18'sd     65;
assign coef[  8] =  18'sd      5;
assign coef[  9] =  18'sd     75;
assign coef[ 10] =  18'sd     94;
assign coef[ 11] =  18'sd     46;
assign coef[ 12] = -18'sd     36;
assign coef[ 13] = -18'sd     94;
assign coef[ 14] = -18'sd     86;
assign coef[ 15] = -18'sd     16;
assign coef[ 16] =  18'sd     67;
assign coef[ 17] =  18'sd    102;
assign coef[ 18] =  18'sd     63;
assign coef[ 19] = -18'sd     23;
assign coef[ 20] = -18'sd     94;
assign coef[ 21] = -18'sd     95;
assign coef[ 22] = -18'sd     25;
assign coef[ 23] =  18'sd     67;
assign coef[ 24] =  18'sd    111;
assign coef[ 25] =  18'sd     71;
assign coef[ 26] = -18'sd     28;
assign coef[ 27] = -18'sd    111;
assign coef[ 28] = -18'sd    115;
assign coef[ 29] = -18'sd     28;
assign coef[ 30] =  18'sd     89;
assign coef[ 31] =  18'sd    149;
assign coef[ 32] =  18'sd    100;
assign coef[ 33] = -18'sd     31;
assign coef[ 34] = -18'sd    152;
assign coef[ 35] = -18'sd    173;
assign coef[ 36] = -18'sd     66;
assign coef[ 37] =  18'sd    101;
assign coef[ 38] =  18'sd    209;
assign coef[ 39] =  18'sd    175;
assign coef[ 40] =  18'sd     11;
assign coef[ 41] = -18'sd    174;
assign coef[ 42] = -18'sd    248;
assign coef[ 43] = -18'sd    150;
assign coef[ 44] =  18'sd     62;
assign coef[ 45] =  18'sd    241;
assign coef[ 46] =  18'sd    257;
assign coef[ 47] =  18'sd     91;
assign coef[ 48] = -18'sd    146;
assign coef[ 49] = -18'sd    286;
assign coef[ 50] = -18'sd    222;
assign coef[ 51] =  18'sd      5;
assign coef[ 52] =  18'sd    234;
assign coef[ 53] =  18'sd    293;
assign coef[ 54] =  18'sd    130;
assign coef[ 55] = -18'sd    140;
assign coef[ 56] = -18'sd    312;
assign coef[ 57] = -18'sd    243;
assign coef[ 58] =  18'sd     33;
assign coef[ 59] =  18'sd    311;
assign coef[ 60] =  18'sd    364;
assign coef[ 61] =  18'sd    115;
assign coef[ 62] = -18'sd    279;
assign coef[ 63] = -18'sd    515;
assign coef[ 64] = -18'sd    370;
assign coef[ 65] =  18'sd    116;
assign coef[ 66] =  18'sd    621;
assign coef[ 67] =  18'sd    745;
assign coef[ 68] =  18'sd    305;
assign coef[ 69] = -18'sd    479;
assign coef[ 70] = -18'sd   1077;
assign coef[ 71] = -18'sd    990;
assign coef[ 72] = -18'sd    136;
assign coef[ 73] =  18'sd   1012;
assign coef[ 74] =  18'sd   1665;
assign coef[ 75] =  18'sd   1240;
assign coef[ 76] = -18'sd    180;
assign coef[ 77] = -18'sd   1772;
assign coef[ 78] = -18'sd   2426;
assign coef[ 79] = -18'sd   1481;
assign coef[ 80] =  18'sd    716;
assign coef[ 81] =  18'sd   2863;
assign coef[ 82] =  18'sd   3433;
assign coef[ 83] =  18'sd   1700;
assign coef[ 84] = -18'sd   1604;
assign coef[ 85] = -18'sd   4499;
assign coef[ 86] = -18'sd   4870;
assign coef[ 87] = -18'sd   1885;
assign coef[ 88] =  18'sd   3161;
assign coef[ 89] =  18'sd   7249;
assign coef[ 90] =  18'sd   7262;
assign coef[ 91] =  18'sd   2026;
assign coef[ 92] = -18'sd   6414;
assign coef[ 93] = -18'sd  13214;
assign coef[ 94] = -18'sd  12866;
assign coef[ 95] = -18'sd   2115;
assign coef[ 96] =  18'sd  17885;
assign coef[ 97] =  18'sd  41412;
assign coef[ 98] =  18'sd  60318;
assign coef[ 99] =  18'sd  67547;
