module ee465_gold_standard_srrc (input sys_clk,
											input sam_clk,
											input [17:0] sig_in,
											output [17:0] sig_out);
											

assign sig_out = sig_in;											

endmodule
