
//RX Filter 18'sd Multiplier Coefficients (headroom)
assign coef[  0] = -18'sd    197;
assign coef[  1] = -18'sd    202;
assign coef[  2] = -18'sd     50;
assign coef[  3] =  18'sd    157;
assign coef[  4] =  18'sd    263;
assign coef[  5] =  18'sd    177;
assign coef[  6] = -18'sd     54;
assign coef[  7] = -18'sd    269;
assign coef[  8] = -18'sd    305;
assign coef[  9] = -18'sd    116;
assign coef[ 10] =  18'sd    178;
assign coef[ 11] =  18'sd    370;
assign coef[ 12] =  18'sd    309;
assign coef[ 13] =  18'sd     19;
assign coef[ 14] = -18'sd    308;
assign coef[ 15] = -18'sd    438;
assign coef[ 16] = -18'sd    264;
assign coef[ 17] =  18'sd    109;
assign coef[ 18] =  18'sd    425;
assign coef[ 19] =  18'sd    454;
assign coef[ 20] =  18'sd    160;
assign coef[ 21] = -18'sd    258;
assign coef[ 22] = -18'sd    504;
assign coef[ 23] = -18'sd    392;
assign coef[ 24] =  18'sd      9;
assign coef[ 25] =  18'sd    413;
assign coef[ 26] =  18'sd    517;
assign coef[ 27] =  18'sd    230;
assign coef[ 28] = -18'sd    247;
assign coef[ 29] = -18'sd    551;
assign coef[ 30] = -18'sd    429;
assign coef[ 31] =  18'sd     57;
assign coef[ 32] =  18'sd    550;
assign coef[ 33] =  18'sd    643;
assign coef[ 34] =  18'sd    203;
assign coef[ 35] = -18'sd    492;
assign coef[ 36] = -18'sd    910;
assign coef[ 37] = -18'sd    654;
assign coef[ 38] =  18'sd    205;
assign coef[ 39] =  18'sd   1098;
assign coef[ 40] =  18'sd   1316;
assign coef[ 41] =  18'sd    539;
assign coef[ 42] = -18'sd    846;
assign coef[ 43] = -18'sd   1902;
assign coef[ 44] = -18'sd   1749;
assign coef[ 45] = -18'sd    241;
assign coef[ 46] =  18'sd   1787;
assign coef[ 47] =  18'sd   2942;
assign coef[ 48] =  18'sd   2190;
assign coef[ 49] = -18'sd    319;
assign coef[ 50] = -18'sd   3131;
assign coef[ 51] = -18'sd   4285;
assign coef[ 52] = -18'sd   2615;
assign coef[ 53] =  18'sd   1265;
assign coef[ 54] =  18'sd   5057;
assign coef[ 55] =  18'sd   6065;
assign coef[ 56] =  18'sd   3003;
assign coef[ 57] = -18'sd   2833;
assign coef[ 58] = -18'sd   7948;
assign coef[ 59] = -18'sd   8603;
assign coef[ 60] = -18'sd   3331;
assign coef[ 61] =  18'sd   5583;
assign coef[ 62] =  18'sd  12805;
assign coef[ 63] =  18'sd  12828;
assign coef[ 64] =  18'sd   3580;
assign coef[ 65] = -18'sd  11331;
assign coef[ 66] = -18'sd  23342;
assign coef[ 67] = -18'sd  22728;
assign coef[ 68] = -18'sd   3735;
assign coef[ 69] =  18'sd  31594;
assign coef[ 70] =  18'sd  73152;
assign coef[ 71] =  18'sd 106550;
assign coef[ 72] =  18'sd 119319;
