
//RX Filter 18'sd Multiplier Coefficients (headroom)
assign coef[  0] =  18'sd      7;
assign coef[  1] = -18'sd     18;
assign coef[  2] = -18'sd     31;
assign coef[  3] = -18'sd     21;
assign coef[  4] =  18'sd      4;
assign coef[  5] =  18'sd     27;
assign coef[  6] =  18'sd     30;
assign coef[  7] =  18'sd     11;
assign coef[  8] = -18'sd     16;
assign coef[  9] = -18'sd     32;
assign coef[ 10] = -18'sd     24;
assign coef[ 11] =  18'sd      2;
assign coef[ 12] =  18'sd     28;
assign coef[ 13] =  18'sd     33;
assign coef[ 14] =  18'sd     14;
assign coef[ 15] = -18'sd     17;
assign coef[ 16] = -18'sd     36;
assign coef[ 17] = -18'sd     29;
assign coef[ 18] =  18'sd      0;
assign coef[ 19] =  18'sd     31;
assign coef[ 20] =  18'sd     40;
assign coef[ 21] =  18'sd     20;
assign coef[ 22] = -18'sd     15;
assign coef[ 23] = -18'sd     41;
assign coef[ 24] = -18'sd     39;
assign coef[ 25] = -18'sd      8;
assign coef[ 26] =  18'sd     30;
assign coef[ 27] =  18'sd     48;
assign coef[ 28] =  18'sd     31;
assign coef[ 29] = -18'sd      8;
assign coef[ 30] = -18'sd     43;
assign coef[ 31] = -18'sd     47;
assign coef[ 32] = -18'sd     18;
assign coef[ 33] =  18'sd     25;
assign coef[ 34] =  18'sd     50;
assign coef[ 35] =  18'sd     40;
assign coef[ 36] =  18'sd      0;
assign coef[ 37] = -18'sd     40;
assign coef[ 38] = -18'sd     51;
assign coef[ 39] = -18'sd     25;
assign coef[ 40] =  18'sd     20;
assign coef[ 41] =  18'sd     51;
assign coef[ 42] =  18'sd     44;
assign coef[ 43] =  18'sd      4;
assign coef[ 44] = -18'sd     40;
assign coef[ 45] = -18'sd     56;
assign coef[ 46] = -18'sd     29;
assign coef[ 47] =  18'sd     21;
assign coef[ 48] =  18'sd     58;
assign coef[ 49] =  18'sd     53;
assign coef[ 50] =  18'sd      7;
assign coef[ 51] = -18'sd     47;
assign coef[ 52] = -18'sd     70;
assign coef[ 53] = -18'sd     42;
assign coef[ 54] =  18'sd     20;
assign coef[ 55] =  18'sd     71;
assign coef[ 56] =  18'sd     73;
assign coef[ 57] =  18'sd     22;
assign coef[ 58] = -18'sd     48;
assign coef[ 59] = -18'sd     87;
assign coef[ 60] = -18'sd     65;
assign coef[ 61] =  18'sd      5;
assign coef[ 62] =  18'sd     75;
assign coef[ 63] =  18'sd     94;
assign coef[ 64] =  18'sd     46;
assign coef[ 65] = -18'sd     36;
assign coef[ 66] = -18'sd     94;
assign coef[ 67] = -18'sd     86;
assign coef[ 68] = -18'sd     16;
assign coef[ 69] =  18'sd     67;
assign coef[ 70] =  18'sd    102;
assign coef[ 71] =  18'sd     63;
assign coef[ 72] = -18'sd     23;
assign coef[ 73] = -18'sd     94;
assign coef[ 74] = -18'sd     95;
assign coef[ 75] = -18'sd     25;
assign coef[ 76] =  18'sd     67;
assign coef[ 77] =  18'sd    111;
assign coef[ 78] =  18'sd     71;
assign coef[ 79] = -18'sd     28;
assign coef[ 80] = -18'sd    111;
assign coef[ 81] = -18'sd    115;
assign coef[ 82] = -18'sd     28;
assign coef[ 83] =  18'sd     89;
assign coef[ 84] =  18'sd    149;
assign coef[ 85] =  18'sd    100;
assign coef[ 86] = -18'sd     31;
assign coef[ 87] = -18'sd    152;
assign coef[ 88] = -18'sd    173;
assign coef[ 89] = -18'sd     66;
assign coef[ 90] =  18'sd    101;
assign coef[ 91] =  18'sd    209;
assign coef[ 92] =  18'sd    175;
assign coef[ 93] =  18'sd     11;
assign coef[ 94] = -18'sd    174;
assign coef[ 95] = -18'sd    248;
assign coef[ 96] = -18'sd    150;
assign coef[ 97] =  18'sd     62;
assign coef[ 98] =  18'sd    241;
assign coef[ 99] =  18'sd    257;
assign coef[100] =  18'sd     91;
assign coef[101] = -18'sd    146;
assign coef[102] = -18'sd    286;
assign coef[103] = -18'sd    222;
assign coef[104] =  18'sd      5;
assign coef[105] =  18'sd    234;
assign coef[106] =  18'sd    293;
assign coef[107] =  18'sd    130;
assign coef[108] = -18'sd    140;
assign coef[109] = -18'sd    312;
assign coef[110] = -18'sd    243;
assign coef[111] =  18'sd     33;
assign coef[112] =  18'sd    311;
assign coef[113] =  18'sd    364;
assign coef[114] =  18'sd    115;
assign coef[115] = -18'sd    279;
assign coef[116] = -18'sd    515;
assign coef[117] = -18'sd    370;
assign coef[118] =  18'sd    116;
assign coef[119] =  18'sd    622;
assign coef[120] =  18'sd    745;
assign coef[121] =  18'sd    305;
assign coef[122] = -18'sd    479;
assign coef[123] = -18'sd   1077;
assign coef[124] = -18'sd    990;
assign coef[125] = -18'sd    136;
assign coef[126] =  18'sd   1012;
assign coef[127] =  18'sd   1666;
assign coef[128] =  18'sd   1240;
assign coef[129] = -18'sd    180;
assign coef[130] = -18'sd   1773;
assign coef[131] = -18'sd   2426;
assign coef[132] = -18'sd   1481;
assign coef[133] =  18'sd    716;
assign coef[134] =  18'sd   2863;
assign coef[135] =  18'sd   3434;
assign coef[136] =  18'sd   1700;
assign coef[137] = -18'sd   1604;
assign coef[138] = -18'sd   4500;
assign coef[139] = -18'sd   4871;
assign coef[140] = -18'sd   1886;
assign coef[141] =  18'sd   3161;
assign coef[142] =  18'sd   7250;
assign coef[143] =  18'sd   7263;
assign coef[144] =  18'sd   2027;
assign coef[145] = -18'sd   6415;
assign coef[146] = -18'sd  13216;
assign coef[147] = -18'sd  12868;
assign coef[148] = -18'sd   2115;
assign coef[149] =  18'sd  17887;
assign coef[150] =  18'sd  41417;
assign coef[151] =  18'sd  60325;
assign coef[152] =  18'sd  67555;
