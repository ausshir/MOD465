
//TX Filter 18'sd Multiplier Coefficients (headroom)
assign coef[  0] =  18'sd     68;
assign coef[  1] =  18'sd    185;
assign coef[  2] =  18'sd    178;
assign coef[  3] =  18'sd     28;
assign coef[  4] = -18'sd    178;
assign coef[  5] = -18'sd    292;
assign coef[  6] = -18'sd    203;
assign coef[  7] =  18'sd     64;
assign coef[  8] =  18'sd    344;
assign coef[  9] =  18'sd    427;
assign coef[ 10] =  18'sd    206;
assign coef[ 11] = -18'sd    220;
assign coef[ 12] = -18'sd    578;
assign coef[ 13] = -18'sd    590;
assign coef[ 14] = -18'sd    173;
assign coef[ 15] =  18'sd    459;
assign coef[ 16] =  18'sd    894;
assign coef[ 17] =  18'sd    778;
assign coef[ 18] =  18'sd     85;
assign coef[ 19] = -18'sd    808;
assign coef[ 20] = -18'sd   1306;
assign coef[ 21] = -18'sd    987;
assign coef[ 22] =  18'sd     82;
assign coef[ 23] =  18'sd   1294;
assign coef[ 24] =  18'sd   1834;
assign coef[ 25] =  18'sd   1209;
assign coef[ 26] = -18'sd    357;
assign coef[ 27] = -18'sd   1957;
assign coef[ 28] = -18'sd   2502;
assign coef[ 29] = -18'sd   1439;
assign coef[ 30] =  18'sd    783;
assign coef[ 31] =  18'sd   2854;
assign coef[ 32] =  18'sd   3348;
assign coef[ 33] =  18'sd   1665;
assign coef[ 34] = -18'sd   1424;
assign coef[ 35] = -18'sd   4079;
assign coef[ 36] = -18'sd   4441;
assign coef[ 37] = -18'sd   1879;
assign coef[ 38] =  18'sd   2390;
assign coef[ 39] =  18'sd   5801;
assign coef[ 40] =  18'sd   5918;
assign coef[ 41] =  18'sd   2071;
assign coef[ 42] = -18'sd   3897;
assign coef[ 43] = -18'sd   8388;
assign coef[ 44] = -18'sd   8096;
assign coef[ 45] = -18'sd   2231;
assign coef[ 46] =  18'sd   6473;
assign coef[ 47] =  18'sd  12798;
assign coef[ 48] =  18'sd  11870;
assign coef[ 49] =  18'sd   2351;
assign coef[ 50] = -18'sd  11844;
assign coef[ 51] = -18'sd  22568;
assign coef[ 52] = -18'sd  21040;
assign coef[ 53] = -18'sd   2426;
assign coef[ 54] =  18'sd  30955;
assign coef[ 55] =  18'sd  69624;
assign coef[ 56] =  18'sd 100453;
assign coef[ 57] =  18'sd 112198;
