
//TX Filter 18'sd P2 LUT Coefficients (headroom)
assign PRECOMP_P2[  0] =  18'sd     68;
assign PRECOMP_P2[  1] =  18'sd    185;
assign PRECOMP_P2[  2] =  18'sd    178;
assign PRECOMP_P2[  3] =  18'sd     28;
assign PRECOMP_P2[  4] = -18'sd    178;
assign PRECOMP_P2[  5] = -18'sd    292;
assign PRECOMP_P2[  6] = -18'sd    203;
assign PRECOMP_P2[  7] =  18'sd     64;
assign PRECOMP_P2[  8] =  18'sd    344;
assign PRECOMP_P2[  9] =  18'sd    427;
assign PRECOMP_P2[ 10] =  18'sd    206;
assign PRECOMP_P2[ 11] = -18'sd    220;
assign PRECOMP_P2[ 12] = -18'sd    578;
assign PRECOMP_P2[ 13] = -18'sd    590;
assign PRECOMP_P2[ 14] = -18'sd    173;
assign PRECOMP_P2[ 15] =  18'sd    459;
assign PRECOMP_P2[ 16] =  18'sd    894;
assign PRECOMP_P2[ 17] =  18'sd    778;
assign PRECOMP_P2[ 18] =  18'sd     85;
assign PRECOMP_P2[ 19] = -18'sd    808;
assign PRECOMP_P2[ 20] = -18'sd   1306;
assign PRECOMP_P2[ 21] = -18'sd    987;
assign PRECOMP_P2[ 22] =  18'sd     82;
assign PRECOMP_P2[ 23] =  18'sd   1294;
assign PRECOMP_P2[ 24] =  18'sd   1834;
assign PRECOMP_P2[ 25] =  18'sd   1209;
assign PRECOMP_P2[ 26] = -18'sd    357;
assign PRECOMP_P2[ 27] = -18'sd   1957;
assign PRECOMP_P2[ 28] = -18'sd   2502;
assign PRECOMP_P2[ 29] = -18'sd   1439;
assign PRECOMP_P2[ 30] =  18'sd    783;
assign PRECOMP_P2[ 31] =  18'sd   2854;
assign PRECOMP_P2[ 32] =  18'sd   3348;
assign PRECOMP_P2[ 33] =  18'sd   1665;
assign PRECOMP_P2[ 34] = -18'sd   1424;
assign PRECOMP_P2[ 35] = -18'sd   4079;
assign PRECOMP_P2[ 36] = -18'sd   4441;
assign PRECOMP_P2[ 37] = -18'sd   1879;
assign PRECOMP_P2[ 38] =  18'sd   2390;
assign PRECOMP_P2[ 39] =  18'sd   5801;
assign PRECOMP_P2[ 40] =  18'sd   5918;
assign PRECOMP_P2[ 41] =  18'sd   2071;
assign PRECOMP_P2[ 42] = -18'sd   3897;
assign PRECOMP_P2[ 43] = -18'sd   8388;
assign PRECOMP_P2[ 44] = -18'sd   8096;
assign PRECOMP_P2[ 45] = -18'sd   2231;
assign PRECOMP_P2[ 46] =  18'sd   6473;
assign PRECOMP_P2[ 47] =  18'sd  12798;
assign PRECOMP_P2[ 48] =  18'sd  11870;
assign PRECOMP_P2[ 49] =  18'sd   2351;
assign PRECOMP_P2[ 50] = -18'sd  11844;
assign PRECOMP_P2[ 51] = -18'sd  22568;
assign PRECOMP_P2[ 52] = -18'sd  21040;
assign PRECOMP_P2[ 53] = -18'sd   2426;
assign PRECOMP_P2[ 54] =  18'sd  30955;
assign PRECOMP_P2[ 55] =  18'sd  69624;
assign PRECOMP_P2[ 56] =  18'sd 100453;
assign PRECOMP_P2[ 57] =  18'sd 112198;
assign PRECOMP_P2[ 58] =  18'sd 100453;
assign PRECOMP_P2[ 59] =  18'sd  69624;
assign PRECOMP_P2[ 60] =  18'sd  30955;
assign PRECOMP_P2[ 61] = -18'sd   2426;
assign PRECOMP_P2[ 62] = -18'sd  21040;
assign PRECOMP_P2[ 63] = -18'sd  22568;
assign PRECOMP_P2[ 64] = -18'sd  11844;
assign PRECOMP_P2[ 65] =  18'sd   2351;
assign PRECOMP_P2[ 66] =  18'sd  11870;
assign PRECOMP_P2[ 67] =  18'sd  12798;
assign PRECOMP_P2[ 68] =  18'sd   6473;
assign PRECOMP_P2[ 69] = -18'sd   2231;
assign PRECOMP_P2[ 70] = -18'sd   8096;
assign PRECOMP_P2[ 71] = -18'sd   8388;
assign PRECOMP_P2[ 72] = -18'sd   3897;
assign PRECOMP_P2[ 73] =  18'sd   2071;
assign PRECOMP_P2[ 74] =  18'sd   5918;
assign PRECOMP_P2[ 75] =  18'sd   5801;
assign PRECOMP_P2[ 76] =  18'sd   2390;
assign PRECOMP_P2[ 77] = -18'sd   1879;
assign PRECOMP_P2[ 78] = -18'sd   4441;
assign PRECOMP_P2[ 79] = -18'sd   4079;
assign PRECOMP_P2[ 80] = -18'sd   1424;
assign PRECOMP_P2[ 81] =  18'sd   1665;
assign PRECOMP_P2[ 82] =  18'sd   3348;
assign PRECOMP_P2[ 83] =  18'sd   2854;
assign PRECOMP_P2[ 84] =  18'sd    783;
assign PRECOMP_P2[ 85] = -18'sd   1439;
assign PRECOMP_P2[ 86] = -18'sd   2502;
assign PRECOMP_P2[ 87] = -18'sd   1957;
assign PRECOMP_P2[ 88] = -18'sd    357;
assign PRECOMP_P2[ 89] =  18'sd   1209;
assign PRECOMP_P2[ 90] =  18'sd   1834;
assign PRECOMP_P2[ 91] =  18'sd   1294;
assign PRECOMP_P2[ 92] =  18'sd     82;
assign PRECOMP_P2[ 93] = -18'sd    987;
assign PRECOMP_P2[ 94] = -18'sd   1306;
assign PRECOMP_P2[ 95] = -18'sd    808;
assign PRECOMP_P2[ 96] =  18'sd     85;
assign PRECOMP_P2[ 97] =  18'sd    778;
assign PRECOMP_P2[ 98] =  18'sd    894;
assign PRECOMP_P2[ 99] =  18'sd    459;
assign PRECOMP_P2[100] = -18'sd    173;
assign PRECOMP_P2[101] = -18'sd    590;
assign PRECOMP_P2[102] = -18'sd    578;
assign PRECOMP_P2[103] = -18'sd    220;
assign PRECOMP_P2[104] =  18'sd    206;
assign PRECOMP_P2[105] =  18'sd    427;
assign PRECOMP_P2[106] =  18'sd    344;
assign PRECOMP_P2[107] =  18'sd     64;
assign PRECOMP_P2[108] = -18'sd    203;
assign PRECOMP_P2[109] = -18'sd    292;
assign PRECOMP_P2[110] = -18'sd    178;
assign PRECOMP_P2[111] =  18'sd     28;
assign PRECOMP_P2[112] =  18'sd    178;
assign PRECOMP_P2[113] =  18'sd    185;
assign PRECOMP_P2[114] =  18'sd     68;



//TX Filter 18'sd P1 LUT Coefficients (headroom)
assign PRECOMP_P1[  0] =  18'sd     46;
assign PRECOMP_P1[  1] =  18'sd    123;
assign PRECOMP_P1[  2] =  18'sd    119;
assign PRECOMP_P1[  3] =  18'sd     19;
assign PRECOMP_P1[  4] = -18'sd    119;
assign PRECOMP_P1[  5] = -18'sd    195;
assign PRECOMP_P1[  6] = -18'sd    136;
assign PRECOMP_P1[  7] =  18'sd     42;
assign PRECOMP_P1[  8] =  18'sd    229;
assign PRECOMP_P1[  9] =  18'sd    285;
assign PRECOMP_P1[ 10] =  18'sd    138;
assign PRECOMP_P1[ 11] = -18'sd    146;
assign PRECOMP_P1[ 12] = -18'sd    385;
assign PRECOMP_P1[ 13] = -18'sd    393;
assign PRECOMP_P1[ 14] = -18'sd    115;
assign PRECOMP_P1[ 15] =  18'sd    306;
assign PRECOMP_P1[ 16] =  18'sd    596;
assign PRECOMP_P1[ 17] =  18'sd    519;
assign PRECOMP_P1[ 18] =  18'sd     56;
assign PRECOMP_P1[ 19] = -18'sd    538;
assign PRECOMP_P1[ 20] = -18'sd    871;
assign PRECOMP_P1[ 21] = -18'sd    658;
assign PRECOMP_P1[ 22] =  18'sd     55;
assign PRECOMP_P1[ 23] =  18'sd    862;
assign PRECOMP_P1[ 24] =  18'sd   1223;
assign PRECOMP_P1[ 25] =  18'sd    806;
assign PRECOMP_P1[ 26] = -18'sd    238;
assign PRECOMP_P1[ 27] = -18'sd   1305;
assign PRECOMP_P1[ 28] = -18'sd   1668;
assign PRECOMP_P1[ 29] = -18'sd    959;
assign PRECOMP_P1[ 30] =  18'sd    522;
assign PRECOMP_P1[ 31] =  18'sd   1903;
assign PRECOMP_P1[ 32] =  18'sd   2232;
assign PRECOMP_P1[ 33] =  18'sd   1110;
assign PRECOMP_P1[ 34] = -18'sd    950;
assign PRECOMP_P1[ 35] = -18'sd   2719;
assign PRECOMP_P1[ 36] = -18'sd   2961;
assign PRECOMP_P1[ 37] = -18'sd   1253;
assign PRECOMP_P1[ 38] =  18'sd   1593;
assign PRECOMP_P1[ 39] =  18'sd   3867;
assign PRECOMP_P1[ 40] =  18'sd   3946;
assign PRECOMP_P1[ 41] =  18'sd   1380;
assign PRECOMP_P1[ 42] = -18'sd   2598;
assign PRECOMP_P1[ 43] = -18'sd   5592;
assign PRECOMP_P1[ 44] = -18'sd   5398;
assign PRECOMP_P1[ 45] = -18'sd   1487;
assign PRECOMP_P1[ 46] =  18'sd   4315;
assign PRECOMP_P1[ 47] =  18'sd   8532;
assign PRECOMP_P1[ 48] =  18'sd   7913;
assign PRECOMP_P1[ 49] =  18'sd   1567;
assign PRECOMP_P1[ 50] = -18'sd   7896;
assign PRECOMP_P1[ 51] = -18'sd  15045;
assign PRECOMP_P1[ 52] = -18'sd  14027;
assign PRECOMP_P1[ 53] = -18'sd   1617;
assign PRECOMP_P1[ 54] =  18'sd  20637;
assign PRECOMP_P1[ 55] =  18'sd  46416;
assign PRECOMP_P1[ 56] =  18'sd  66969;
assign PRECOMP_P1[ 57] =  18'sd  74799;
assign PRECOMP_P1[ 58] =  18'sd  66969;
assign PRECOMP_P1[ 59] =  18'sd  46416;
assign PRECOMP_P1[ 60] =  18'sd  20637;
assign PRECOMP_P1[ 61] = -18'sd   1617;
assign PRECOMP_P1[ 62] = -18'sd  14027;
assign PRECOMP_P1[ 63] = -18'sd  15045;
assign PRECOMP_P1[ 64] = -18'sd   7896;
assign PRECOMP_P1[ 65] =  18'sd   1567;
assign PRECOMP_P1[ 66] =  18'sd   7913;
assign PRECOMP_P1[ 67] =  18'sd   8532;
assign PRECOMP_P1[ 68] =  18'sd   4315;
assign PRECOMP_P1[ 69] = -18'sd   1487;
assign PRECOMP_P1[ 70] = -18'sd   5398;
assign PRECOMP_P1[ 71] = -18'sd   5592;
assign PRECOMP_P1[ 72] = -18'sd   2598;
assign PRECOMP_P1[ 73] =  18'sd   1380;
assign PRECOMP_P1[ 74] =  18'sd   3946;
assign PRECOMP_P1[ 75] =  18'sd   3867;
assign PRECOMP_P1[ 76] =  18'sd   1593;
assign PRECOMP_P1[ 77] = -18'sd   1253;
assign PRECOMP_P1[ 78] = -18'sd   2961;
assign PRECOMP_P1[ 79] = -18'sd   2719;
assign PRECOMP_P1[ 80] = -18'sd    950;
assign PRECOMP_P1[ 81] =  18'sd   1110;
assign PRECOMP_P1[ 82] =  18'sd   2232;
assign PRECOMP_P1[ 83] =  18'sd   1903;
assign PRECOMP_P1[ 84] =  18'sd    522;
assign PRECOMP_P1[ 85] = -18'sd    959;
assign PRECOMP_P1[ 86] = -18'sd   1668;
assign PRECOMP_P1[ 87] = -18'sd   1305;
assign PRECOMP_P1[ 88] = -18'sd    238;
assign PRECOMP_P1[ 89] =  18'sd    806;
assign PRECOMP_P1[ 90] =  18'sd   1223;
assign PRECOMP_P1[ 91] =  18'sd    862;
assign PRECOMP_P1[ 92] =  18'sd     55;
assign PRECOMP_P1[ 93] = -18'sd    658;
assign PRECOMP_P1[ 94] = -18'sd    871;
assign PRECOMP_P1[ 95] = -18'sd    538;
assign PRECOMP_P1[ 96] =  18'sd     56;
assign PRECOMP_P1[ 97] =  18'sd    519;
assign PRECOMP_P1[ 98] =  18'sd    596;
assign PRECOMP_P1[ 99] =  18'sd    306;
assign PRECOMP_P1[100] = -18'sd    115;
assign PRECOMP_P1[101] = -18'sd    393;
assign PRECOMP_P1[102] = -18'sd    385;
assign PRECOMP_P1[103] = -18'sd    146;
assign PRECOMP_P1[104] =  18'sd    138;
assign PRECOMP_P1[105] =  18'sd    285;
assign PRECOMP_P1[106] =  18'sd    229;
assign PRECOMP_P1[107] =  18'sd     42;
assign PRECOMP_P1[108] = -18'sd    136;
assign PRECOMP_P1[109] = -18'sd    195;
assign PRECOMP_P1[110] = -18'sd    119;
assign PRECOMP_P1[111] =  18'sd     19;
assign PRECOMP_P1[112] =  18'sd    119;
assign PRECOMP_P1[113] =  18'sd    123;
assign PRECOMP_P1[114] =  18'sd     46;



//TX Filter 18'sd N1 LUT Coefficients (headroom)
assign PRECOMP_N1[  0] = -18'sd     46;
assign PRECOMP_N1[  1] = -18'sd    123;
assign PRECOMP_N1[  2] = -18'sd    119;
assign PRECOMP_N1[  3] = -18'sd     19;
assign PRECOMP_N1[  4] =  18'sd    119;
assign PRECOMP_N1[  5] =  18'sd    195;
assign PRECOMP_N1[  6] =  18'sd    136;
assign PRECOMP_N1[  7] = -18'sd     42;
assign PRECOMP_N1[  8] = -18'sd    229;
assign PRECOMP_N1[  9] = -18'sd    285;
assign PRECOMP_N1[ 10] = -18'sd    138;
assign PRECOMP_N1[ 11] =  18'sd    146;
assign PRECOMP_N1[ 12] =  18'sd    385;
assign PRECOMP_N1[ 13] =  18'sd    393;
assign PRECOMP_N1[ 14] =  18'sd    115;
assign PRECOMP_N1[ 15] = -18'sd    306;
assign PRECOMP_N1[ 16] = -18'sd    596;
assign PRECOMP_N1[ 17] = -18'sd    519;
assign PRECOMP_N1[ 18] = -18'sd     56;
assign PRECOMP_N1[ 19] =  18'sd    538;
assign PRECOMP_N1[ 20] =  18'sd    871;
assign PRECOMP_N1[ 21] =  18'sd    658;
assign PRECOMP_N1[ 22] = -18'sd     55;
assign PRECOMP_N1[ 23] = -18'sd    862;
assign PRECOMP_N1[ 24] = -18'sd   1223;
assign PRECOMP_N1[ 25] = -18'sd    806;
assign PRECOMP_N1[ 26] =  18'sd    238;
assign PRECOMP_N1[ 27] =  18'sd   1305;
assign PRECOMP_N1[ 28] =  18'sd   1668;
assign PRECOMP_N1[ 29] =  18'sd    959;
assign PRECOMP_N1[ 30] = -18'sd    522;
assign PRECOMP_N1[ 31] = -18'sd   1903;
assign PRECOMP_N1[ 32] = -18'sd   2232;
assign PRECOMP_N1[ 33] = -18'sd   1110;
assign PRECOMP_N1[ 34] =  18'sd    950;
assign PRECOMP_N1[ 35] =  18'sd   2719;
assign PRECOMP_N1[ 36] =  18'sd   2961;
assign PRECOMP_N1[ 37] =  18'sd   1253;
assign PRECOMP_N1[ 38] = -18'sd   1593;
assign PRECOMP_N1[ 39] = -18'sd   3867;
assign PRECOMP_N1[ 40] = -18'sd   3946;
assign PRECOMP_N1[ 41] = -18'sd   1380;
assign PRECOMP_N1[ 42] =  18'sd   2598;
assign PRECOMP_N1[ 43] =  18'sd   5592;
assign PRECOMP_N1[ 44] =  18'sd   5398;
assign PRECOMP_N1[ 45] =  18'sd   1487;
assign PRECOMP_N1[ 46] = -18'sd   4315;
assign PRECOMP_N1[ 47] = -18'sd   8532;
assign PRECOMP_N1[ 48] = -18'sd   7913;
assign PRECOMP_N1[ 49] = -18'sd   1567;
assign PRECOMP_N1[ 50] =  18'sd   7896;
assign PRECOMP_N1[ 51] =  18'sd  15045;
assign PRECOMP_N1[ 52] =  18'sd  14027;
assign PRECOMP_N1[ 53] =  18'sd   1617;
assign PRECOMP_N1[ 54] = -18'sd  20637;
assign PRECOMP_N1[ 55] = -18'sd  46416;
assign PRECOMP_N1[ 56] = -18'sd  66969;
assign PRECOMP_N1[ 57] = -18'sd  74799;
assign PRECOMP_N1[ 58] = -18'sd  66969;
assign PRECOMP_N1[ 59] = -18'sd  46416;
assign PRECOMP_N1[ 60] = -18'sd  20637;
assign PRECOMP_N1[ 61] =  18'sd   1617;
assign PRECOMP_N1[ 62] =  18'sd  14027;
assign PRECOMP_N1[ 63] =  18'sd  15045;
assign PRECOMP_N1[ 64] =  18'sd   7896;
assign PRECOMP_N1[ 65] = -18'sd   1567;
assign PRECOMP_N1[ 66] = -18'sd   7913;
assign PRECOMP_N1[ 67] = -18'sd   8532;
assign PRECOMP_N1[ 68] = -18'sd   4315;
assign PRECOMP_N1[ 69] =  18'sd   1487;
assign PRECOMP_N1[ 70] =  18'sd   5398;
assign PRECOMP_N1[ 71] =  18'sd   5592;
assign PRECOMP_N1[ 72] =  18'sd   2598;
assign PRECOMP_N1[ 73] = -18'sd   1380;
assign PRECOMP_N1[ 74] = -18'sd   3946;
assign PRECOMP_N1[ 75] = -18'sd   3867;
assign PRECOMP_N1[ 76] = -18'sd   1593;
assign PRECOMP_N1[ 77] =  18'sd   1253;
assign PRECOMP_N1[ 78] =  18'sd   2961;
assign PRECOMP_N1[ 79] =  18'sd   2719;
assign PRECOMP_N1[ 80] =  18'sd    950;
assign PRECOMP_N1[ 81] = -18'sd   1110;
assign PRECOMP_N1[ 82] = -18'sd   2232;
assign PRECOMP_N1[ 83] = -18'sd   1903;
assign PRECOMP_N1[ 84] = -18'sd    522;
assign PRECOMP_N1[ 85] =  18'sd    959;
assign PRECOMP_N1[ 86] =  18'sd   1668;
assign PRECOMP_N1[ 87] =  18'sd   1305;
assign PRECOMP_N1[ 88] =  18'sd    238;
assign PRECOMP_N1[ 89] = -18'sd    806;
assign PRECOMP_N1[ 90] = -18'sd   1223;
assign PRECOMP_N1[ 91] = -18'sd    862;
assign PRECOMP_N1[ 92] = -18'sd     55;
assign PRECOMP_N1[ 93] =  18'sd    658;
assign PRECOMP_N1[ 94] =  18'sd    871;
assign PRECOMP_N1[ 95] =  18'sd    538;
assign PRECOMP_N1[ 96] = -18'sd     56;
assign PRECOMP_N1[ 97] = -18'sd    519;
assign PRECOMP_N1[ 98] = -18'sd    596;
assign PRECOMP_N1[ 99] = -18'sd    306;
assign PRECOMP_N1[100] =  18'sd    115;
assign PRECOMP_N1[101] =  18'sd    393;
assign PRECOMP_N1[102] =  18'sd    385;
assign PRECOMP_N1[103] =  18'sd    146;
assign PRECOMP_N1[104] = -18'sd    138;
assign PRECOMP_N1[105] = -18'sd    285;
assign PRECOMP_N1[106] = -18'sd    229;
assign PRECOMP_N1[107] = -18'sd     42;
assign PRECOMP_N1[108] =  18'sd    136;
assign PRECOMP_N1[109] =  18'sd    195;
assign PRECOMP_N1[110] =  18'sd    119;
assign PRECOMP_N1[111] = -18'sd     19;
assign PRECOMP_N1[112] = -18'sd    119;
assign PRECOMP_N1[113] = -18'sd    123;
assign PRECOMP_N1[114] = -18'sd     46;



//TX Filter 18'sd N2 LUT Coefficients (headroom)
assign PRECOMP_N2[  0] = -18'sd     68;
assign PRECOMP_N2[  1] = -18'sd    185;
assign PRECOMP_N2[  2] = -18'sd    178;
assign PRECOMP_N2[  3] = -18'sd     28;
assign PRECOMP_N2[  4] =  18'sd    178;
assign PRECOMP_N2[  5] =  18'sd    292;
assign PRECOMP_N2[  6] =  18'sd    203;
assign PRECOMP_N2[  7] = -18'sd     64;
assign PRECOMP_N2[  8] = -18'sd    344;
assign PRECOMP_N2[  9] = -18'sd    427;
assign PRECOMP_N2[ 10] = -18'sd    206;
assign PRECOMP_N2[ 11] =  18'sd    220;
assign PRECOMP_N2[ 12] =  18'sd    578;
assign PRECOMP_N2[ 13] =  18'sd    590;
assign PRECOMP_N2[ 14] =  18'sd    173;
assign PRECOMP_N2[ 15] = -18'sd    459;
assign PRECOMP_N2[ 16] = -18'sd    894;
assign PRECOMP_N2[ 17] = -18'sd    778;
assign PRECOMP_N2[ 18] = -18'sd     85;
assign PRECOMP_N2[ 19] =  18'sd    808;
assign PRECOMP_N2[ 20] =  18'sd   1306;
assign PRECOMP_N2[ 21] =  18'sd    987;
assign PRECOMP_N2[ 22] = -18'sd     82;
assign PRECOMP_N2[ 23] = -18'sd   1294;
assign PRECOMP_N2[ 24] = -18'sd   1834;
assign PRECOMP_N2[ 25] = -18'sd   1209;
assign PRECOMP_N2[ 26] =  18'sd    357;
assign PRECOMP_N2[ 27] =  18'sd   1957;
assign PRECOMP_N2[ 28] =  18'sd   2502;
assign PRECOMP_N2[ 29] =  18'sd   1439;
assign PRECOMP_N2[ 30] = -18'sd    783;
assign PRECOMP_N2[ 31] = -18'sd   2854;
assign PRECOMP_N2[ 32] = -18'sd   3348;
assign PRECOMP_N2[ 33] = -18'sd   1665;
assign PRECOMP_N2[ 34] =  18'sd   1424;
assign PRECOMP_N2[ 35] =  18'sd   4079;
assign PRECOMP_N2[ 36] =  18'sd   4441;
assign PRECOMP_N2[ 37] =  18'sd   1879;
assign PRECOMP_N2[ 38] = -18'sd   2390;
assign PRECOMP_N2[ 39] = -18'sd   5801;
assign PRECOMP_N2[ 40] = -18'sd   5918;
assign PRECOMP_N2[ 41] = -18'sd   2071;
assign PRECOMP_N2[ 42] =  18'sd   3897;
assign PRECOMP_N2[ 43] =  18'sd   8388;
assign PRECOMP_N2[ 44] =  18'sd   8096;
assign PRECOMP_N2[ 45] =  18'sd   2231;
assign PRECOMP_N2[ 46] = -18'sd   6473;
assign PRECOMP_N2[ 47] = -18'sd  12798;
assign PRECOMP_N2[ 48] = -18'sd  11870;
assign PRECOMP_N2[ 49] = -18'sd   2351;
assign PRECOMP_N2[ 50] =  18'sd  11844;
assign PRECOMP_N2[ 51] =  18'sd  22568;
assign PRECOMP_N2[ 52] =  18'sd  21040;
assign PRECOMP_N2[ 53] =  18'sd   2426;
assign PRECOMP_N2[ 54] = -18'sd  30955;
assign PRECOMP_N2[ 55] = -18'sd  69624;
assign PRECOMP_N2[ 56] = -18'sd 100453;
assign PRECOMP_N2[ 57] = -18'sd 112198;
assign PRECOMP_N2[ 58] = -18'sd 100453;
assign PRECOMP_N2[ 59] = -18'sd  69624;
assign PRECOMP_N2[ 60] = -18'sd  30955;
assign PRECOMP_N2[ 61] =  18'sd   2426;
assign PRECOMP_N2[ 62] =  18'sd  21040;
assign PRECOMP_N2[ 63] =  18'sd  22568;
assign PRECOMP_N2[ 64] =  18'sd  11844;
assign PRECOMP_N2[ 65] = -18'sd   2351;
assign PRECOMP_N2[ 66] = -18'sd  11870;
assign PRECOMP_N2[ 67] = -18'sd  12798;
assign PRECOMP_N2[ 68] = -18'sd   6473;
assign PRECOMP_N2[ 69] =  18'sd   2231;
assign PRECOMP_N2[ 70] =  18'sd   8096;
assign PRECOMP_N2[ 71] =  18'sd   8388;
assign PRECOMP_N2[ 72] =  18'sd   3897;
assign PRECOMP_N2[ 73] = -18'sd   2071;
assign PRECOMP_N2[ 74] = -18'sd   5918;
assign PRECOMP_N2[ 75] = -18'sd   5801;
assign PRECOMP_N2[ 76] = -18'sd   2390;
assign PRECOMP_N2[ 77] =  18'sd   1879;
assign PRECOMP_N2[ 78] =  18'sd   4441;
assign PRECOMP_N2[ 79] =  18'sd   4079;
assign PRECOMP_N2[ 80] =  18'sd   1424;
assign PRECOMP_N2[ 81] = -18'sd   1665;
assign PRECOMP_N2[ 82] = -18'sd   3348;
assign PRECOMP_N2[ 83] = -18'sd   2854;
assign PRECOMP_N2[ 84] = -18'sd    783;
assign PRECOMP_N2[ 85] =  18'sd   1439;
assign PRECOMP_N2[ 86] =  18'sd   2502;
assign PRECOMP_N2[ 87] =  18'sd   1957;
assign PRECOMP_N2[ 88] =  18'sd    357;
assign PRECOMP_N2[ 89] = -18'sd   1209;
assign PRECOMP_N2[ 90] = -18'sd   1834;
assign PRECOMP_N2[ 91] = -18'sd   1294;
assign PRECOMP_N2[ 92] = -18'sd     82;
assign PRECOMP_N2[ 93] =  18'sd    987;
assign PRECOMP_N2[ 94] =  18'sd   1306;
assign PRECOMP_N2[ 95] =  18'sd    808;
assign PRECOMP_N2[ 96] = -18'sd     85;
assign PRECOMP_N2[ 97] = -18'sd    778;
assign PRECOMP_N2[ 98] = -18'sd    894;
assign PRECOMP_N2[ 99] = -18'sd    459;
assign PRECOMP_N2[100] =  18'sd    173;
assign PRECOMP_N2[101] =  18'sd    590;
assign PRECOMP_N2[102] =  18'sd    578;
assign PRECOMP_N2[103] =  18'sd    220;
assign PRECOMP_N2[104] = -18'sd    206;
assign PRECOMP_N2[105] = -18'sd    427;
assign PRECOMP_N2[106] = -18'sd    344;
assign PRECOMP_N2[107] = -18'sd     64;
assign PRECOMP_N2[108] =  18'sd    203;
assign PRECOMP_N2[109] =  18'sd    292;
assign PRECOMP_N2[110] =  18'sd    178;
assign PRECOMP_N2[111] = -18'sd     28;
assign PRECOMP_N2[112] = -18'sd    178;
assign PRECOMP_N2[113] = -18'sd    185;
assign PRECOMP_N2[114] = -18'sd     68;

