
//TX Filter 18'sd Multiplier Coefficients (headroom)
assign coef[  0] = -18'sd     59;
assign coef[  1] = -18'sd     19;
assign coef[  2] =  18'sd     49;
assign coef[  3] =  18'sd    102;
assign coef[  4] =  18'sd     96;
assign coef[  5] =  18'sd     17;
assign coef[  6] = -18'sd     97;
assign coef[  7] = -18'sd    174;
assign coef[  8] = -18'sd    145;
assign coef[  9] = -18'sd      5;
assign coef[ 10] =  18'sd    174;
assign coef[ 11] =  18'sd    274;
assign coef[ 12] =  18'sd    206;
assign coef[ 13] = -18'sd     23;
assign coef[ 14] = -18'sd    287;
assign coef[ 15] = -18'sd    411;
assign coef[ 16] = -18'sd    277;
assign coef[ 17] =  18'sd     75;
assign coef[ 18] =  18'sd    448;
assign coef[ 19] =  18'sd    590;
assign coef[ 20] =  18'sd    359;
assign coef[ 21] = -18'sd    160;
assign coef[ 22] = -18'sd    669;
assign coef[ 23] = -18'sd    821;
assign coef[ 24] = -18'sd    449;
assign coef[ 25] =  18'sd    291;
assign coef[ 26] =  18'sd    966;
assign coef[ 27] =  18'sd   1114;
assign coef[ 28] =  18'sd    545;
assign coef[ 29] = -18'sd    484;
assign coef[ 30] = -18'sd   1363;
assign coef[ 31] = -18'sd   1485;
assign coef[ 32] = -18'sd    643;
assign coef[ 33] =  18'sd    762;
assign coef[ 34] =  18'sd   1893;
assign coef[ 35] =  18'sd   1956;
assign coef[ 36] =  18'sd    739;
assign coef[ 37] = -18'sd   1164;
assign coef[ 38] = -18'sd   2609;
assign coef[ 39] = -18'sd   2571;
assign coef[ 40] = -18'sd    830;
assign coef[ 41] =  18'sd   1751;
assign coef[ 42] =  18'sd   3616;
assign coef[ 43] =  18'sd   3412;
assign coef[ 44] =  18'sd    911;
assign coef[ 45] = -18'sd   2654;
assign coef[ 46] = -18'sd   5130;
assign coef[ 47] = -18'sd   4669;
assign coef[ 48] = -18'sd    979;
assign coef[ 49] =  18'sd   4186;
assign coef[ 50] =  18'sd   7726;
assign coef[ 51] =  18'sd   6878;
assign coef[ 52] =  18'sd   1030;
assign coef[ 53] = -18'sd   7375;
assign coef[ 54] = -18'sd  13512;
assign coef[ 55] = -18'sd  12306;
assign coef[ 56] = -18'sd   1062;
assign coef[ 57] =  18'sd  18745;
assign coef[ 58] =  18'sd  41517;
assign coef[ 59] =  18'sd  59604;
assign coef[ 60] =  18'sd  66483;
