
//TX Filter 18'sd Multiplier Coefficients (headroom)
assign coef[  0] = -18'sd    115;
assign coef[  1] = -18'sd    152;
assign coef[  2] = -18'sd     74;
assign coef[  3] =  18'sd     78;
assign coef[  4] =  18'sd    199;
assign coef[  5] =  18'sd    186;
assign coef[  6] =  18'sd     24;
assign coef[  7] = -18'sd    193;
assign coef[  8] = -18'sd    308;
assign coef[  9] = -18'sd    209;
assign coef[ 10] =  18'sd     74;
assign coef[ 11] =  18'sd    364;
assign coef[ 12] =  18'sd    445;
assign coef[ 13] =  18'sd    209;
assign coef[ 14] = -18'sd    235;
assign coef[ 15] = -18'sd    603;
assign coef[ 16] = -18'sd    608;
assign coef[ 17] = -18'sd    171;
assign coef[ 18] =  18'sd    481;
assign coef[ 19] =  18'sd    922;
assign coef[ 20] =  18'sd    795;
assign coef[ 21] =  18'sd     79;
assign coef[ 22] = -18'sd    834;
assign coef[ 23] = -18'sd   1337;
assign coef[ 24] = -18'sd   1001;
assign coef[ 25] =  18'sd     93;
assign coef[ 26] =  18'sd   1323;
assign coef[ 27] =  18'sd   1864;
assign coef[ 28] =  18'sd   1221;
assign coef[ 29] = -18'sd    372;
assign coef[ 30] = -18'sd   1988;
assign coef[ 31] = -18'sd   2529;
assign coef[ 32] = -18'sd   1446;
assign coef[ 33] =  18'sd    801;
assign coef[ 34] =  18'sd   2884;
assign coef[ 35] =  18'sd   3370;
assign coef[ 36] =  18'sd   1667;
assign coef[ 37] = -18'sd   1443;
assign coef[ 38] = -18'sd   4104;
assign coef[ 39] = -18'sd   4456;
assign coef[ 40] = -18'sd   1875;
assign coef[ 41] =  18'sd   2407;
assign coef[ 42] =  18'sd   5818;
assign coef[ 43] =  18'sd   5923;
assign coef[ 44] =  18'sd   2061;
assign coef[ 45] = -18'sd   3910;
assign coef[ 46] = -18'sd   8392;
assign coef[ 47] = -18'sd   8087;
assign coef[ 48] = -18'sd   2217;
assign coef[ 49] =  18'sd   6477;
assign coef[ 50] =  18'sd  12782;
assign coef[ 51] =  18'sd  11841;
assign coef[ 52] =  18'sd   2333;
assign coef[ 53] = -18'sd  11827;
assign coef[ 54] = -18'sd  22513;
assign coef[ 55] = -18'sd  20976;
assign coef[ 56] = -18'sd   2406;
assign coef[ 57] =  18'sd  30874;
assign coef[ 58] =  18'sd  69414;
assign coef[ 59] =  18'sd 100135;
assign coef[ 60] =  18'sd 111838;
