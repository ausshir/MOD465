
//TX Filter 18'sd P2 LUT Coefficients (headroom)
assign PRECOMP_P2[  0] = -18'sd     29;
assign PRECOMP_P2[  1] = -18'sd     10;
assign PRECOMP_P2[  2] =  18'sd     24;
assign PRECOMP_P2[  3] =  18'sd     51;
assign PRECOMP_P2[  4] =  18'sd     48;
assign PRECOMP_P2[  5] =  18'sd      9;
assign PRECOMP_P2[  6] = -18'sd     49;
assign PRECOMP_P2[  7] = -18'sd     87;
assign PRECOMP_P2[  8] = -18'sd     73;
assign PRECOMP_P2[  9] = -18'sd      3;
assign PRECOMP_P2[ 10] =  18'sd     87;
assign PRECOMP_P2[ 11] =  18'sd    137;
assign PRECOMP_P2[ 12] =  18'sd    103;
assign PRECOMP_P2[ 13] = -18'sd     11;
assign PRECOMP_P2[ 14] = -18'sd    144;
assign PRECOMP_P2[ 15] = -18'sd    205;
assign PRECOMP_P2[ 16] = -18'sd    139;
assign PRECOMP_P2[ 17] =  18'sd     37;
assign PRECOMP_P2[ 18] =  18'sd    224;
assign PRECOMP_P2[ 19] =  18'sd    295;
assign PRECOMP_P2[ 20] =  18'sd    180;
assign PRECOMP_P2[ 21] = -18'sd     80;
assign PRECOMP_P2[ 22] = -18'sd    334;
assign PRECOMP_P2[ 23] = -18'sd    410;
assign PRECOMP_P2[ 24] = -18'sd    225;
assign PRECOMP_P2[ 25] =  18'sd    145;
assign PRECOMP_P2[ 26] =  18'sd    483;
assign PRECOMP_P2[ 27] =  18'sd    557;
assign PRECOMP_P2[ 28] =  18'sd    272;
assign PRECOMP_P2[ 29] = -18'sd    242;
assign PRECOMP_P2[ 30] = -18'sd    682;
assign PRECOMP_P2[ 31] = -18'sd    742;
assign PRECOMP_P2[ 32] = -18'sd    321;
assign PRECOMP_P2[ 33] =  18'sd    381;
assign PRECOMP_P2[ 34] =  18'sd    946;
assign PRECOMP_P2[ 35] =  18'sd    978;
assign PRECOMP_P2[ 36] =  18'sd    370;
assign PRECOMP_P2[ 37] = -18'sd    582;
assign PRECOMP_P2[ 38] = -18'sd   1305;
assign PRECOMP_P2[ 39] = -18'sd   1286;
assign PRECOMP_P2[ 40] = -18'sd    415;
assign PRECOMP_P2[ 41] =  18'sd    876;
assign PRECOMP_P2[ 42] =  18'sd   1808;
assign PRECOMP_P2[ 43] =  18'sd   1706;
assign PRECOMP_P2[ 44] =  18'sd    456;
assign PRECOMP_P2[ 45] = -18'sd   1327;
assign PRECOMP_P2[ 46] = -18'sd   2565;
assign PRECOMP_P2[ 47] = -18'sd   2335;
assign PRECOMP_P2[ 48] = -18'sd    490;
assign PRECOMP_P2[ 49] =  18'sd   2093;
assign PRECOMP_P2[ 50] =  18'sd   3863;
assign PRECOMP_P2[ 51] =  18'sd   3439;
assign PRECOMP_P2[ 52] =  18'sd    515;
assign PRECOMP_P2[ 53] = -18'sd   3687;
assign PRECOMP_P2[ 54] = -18'sd   6756;
assign PRECOMP_P2[ 55] = -18'sd   6153;
assign PRECOMP_P2[ 56] = -18'sd    531;
assign PRECOMP_P2[ 57] =  18'sd   9372;
assign PRECOMP_P2[ 58] =  18'sd  20759;
assign PRECOMP_P2[ 59] =  18'sd  29802;
assign PRECOMP_P2[ 60] =  18'sd  33241;
assign PRECOMP_P2[ 61] =  18'sd  29802;
assign PRECOMP_P2[ 62] =  18'sd  20759;
assign PRECOMP_P2[ 63] =  18'sd   9372;
assign PRECOMP_P2[ 64] = -18'sd    531;
assign PRECOMP_P2[ 65] = -18'sd   6153;
assign PRECOMP_P2[ 66] = -18'sd   6756;
assign PRECOMP_P2[ 67] = -18'sd   3687;
assign PRECOMP_P2[ 68] =  18'sd    515;
assign PRECOMP_P2[ 69] =  18'sd   3439;
assign PRECOMP_P2[ 70] =  18'sd   3863;
assign PRECOMP_P2[ 71] =  18'sd   2093;
assign PRECOMP_P2[ 72] = -18'sd    490;
assign PRECOMP_P2[ 73] = -18'sd   2335;
assign PRECOMP_P2[ 74] = -18'sd   2565;
assign PRECOMP_P2[ 75] = -18'sd   1327;
assign PRECOMP_P2[ 76] =  18'sd    456;
assign PRECOMP_P2[ 77] =  18'sd   1706;
assign PRECOMP_P2[ 78] =  18'sd   1808;
assign PRECOMP_P2[ 79] =  18'sd    876;
assign PRECOMP_P2[ 80] = -18'sd    415;
assign PRECOMP_P2[ 81] = -18'sd   1286;
assign PRECOMP_P2[ 82] = -18'sd   1305;
assign PRECOMP_P2[ 83] = -18'sd    582;
assign PRECOMP_P2[ 84] =  18'sd    370;
assign PRECOMP_P2[ 85] =  18'sd    978;
assign PRECOMP_P2[ 86] =  18'sd    946;
assign PRECOMP_P2[ 87] =  18'sd    381;
assign PRECOMP_P2[ 88] = -18'sd    321;
assign PRECOMP_P2[ 89] = -18'sd    742;
assign PRECOMP_P2[ 90] = -18'sd    682;
assign PRECOMP_P2[ 91] = -18'sd    242;
assign PRECOMP_P2[ 92] =  18'sd    272;
assign PRECOMP_P2[ 93] =  18'sd    557;
assign PRECOMP_P2[ 94] =  18'sd    483;
assign PRECOMP_P2[ 95] =  18'sd    145;
assign PRECOMP_P2[ 96] = -18'sd    225;
assign PRECOMP_P2[ 97] = -18'sd    410;
assign PRECOMP_P2[ 98] = -18'sd    334;
assign PRECOMP_P2[ 99] = -18'sd     80;
assign PRECOMP_P2[100] =  18'sd    180;
assign PRECOMP_P2[101] =  18'sd    295;
assign PRECOMP_P2[102] =  18'sd    224;
assign PRECOMP_P2[103] =  18'sd     37;
assign PRECOMP_P2[104] = -18'sd    139;
assign PRECOMP_P2[105] = -18'sd    205;
assign PRECOMP_P2[106] = -18'sd    144;
assign PRECOMP_P2[107] = -18'sd     11;
assign PRECOMP_P2[108] =  18'sd    103;
assign PRECOMP_P2[109] =  18'sd    137;
assign PRECOMP_P2[110] =  18'sd     87;
assign PRECOMP_P2[111] = -18'sd      3;
assign PRECOMP_P2[112] = -18'sd     73;
assign PRECOMP_P2[113] = -18'sd     87;
assign PRECOMP_P2[114] = -18'sd     49;
assign PRECOMP_P2[115] =  18'sd      9;
assign PRECOMP_P2[116] =  18'sd     48;
assign PRECOMP_P2[117] =  18'sd     51;
assign PRECOMP_P2[118] =  18'sd     24;
assign PRECOMP_P2[119] = -18'sd     10;
assign PRECOMP_P2[120] = -18'sd     29;



//TX Filter 18'sd P1 LUT Coefficients (headroom)
assign PRECOMP_P1[  0] = -18'sd     10;
assign PRECOMP_P1[  1] = -18'sd      3;
assign PRECOMP_P1[  2] =  18'sd      8;
assign PRECOMP_P1[  3] =  18'sd     17;
assign PRECOMP_P1[  4] =  18'sd     16;
assign PRECOMP_P1[  5] =  18'sd      3;
assign PRECOMP_P1[  6] = -18'sd     16;
assign PRECOMP_P1[  7] = -18'sd     29;
assign PRECOMP_P1[  8] = -18'sd     24;
assign PRECOMP_P1[  9] = -18'sd      1;
assign PRECOMP_P1[ 10] =  18'sd     29;
assign PRECOMP_P1[ 11] =  18'sd     46;
assign PRECOMP_P1[ 12] =  18'sd     34;
assign PRECOMP_P1[ 13] = -18'sd      4;
assign PRECOMP_P1[ 14] = -18'sd     48;
assign PRECOMP_P1[ 15] = -18'sd     69;
assign PRECOMP_P1[ 16] = -18'sd     46;
assign PRECOMP_P1[ 17] =  18'sd     12;
assign PRECOMP_P1[ 18] =  18'sd     75;
assign PRECOMP_P1[ 19] =  18'sd     99;
assign PRECOMP_P1[ 20] =  18'sd     60;
assign PRECOMP_P1[ 21] = -18'sd     27;
assign PRECOMP_P1[ 22] = -18'sd    112;
assign PRECOMP_P1[ 23] = -18'sd    137;
assign PRECOMP_P1[ 24] = -18'sd     75;
assign PRECOMP_P1[ 25] =  18'sd     49;
assign PRECOMP_P1[ 26] =  18'sd    161;
assign PRECOMP_P1[ 27] =  18'sd    186;
assign PRECOMP_P1[ 28] =  18'sd     91;
assign PRECOMP_P1[ 29] = -18'sd     81;
assign PRECOMP_P1[ 30] = -18'sd    228;
assign PRECOMP_P1[ 31] = -18'sd    248;
assign PRECOMP_P1[ 32] = -18'sd    107;
assign PRECOMP_P1[ 33] =  18'sd    127;
assign PRECOMP_P1[ 34] =  18'sd    316;
assign PRECOMP_P1[ 35] =  18'sd    327;
assign PRECOMP_P1[ 36] =  18'sd    123;
assign PRECOMP_P1[ 37] = -18'sd    194;
assign PRECOMP_P1[ 38] = -18'sd    436;
assign PRECOMP_P1[ 39] = -18'sd    429;
assign PRECOMP_P1[ 40] = -18'sd    139;
assign PRECOMP_P1[ 41] =  18'sd    292;
assign PRECOMP_P1[ 42] =  18'sd    604;
assign PRECOMP_P1[ 43] =  18'sd    570;
assign PRECOMP_P1[ 44] =  18'sd    152;
assign PRECOMP_P1[ 45] = -18'sd    443;
assign PRECOMP_P1[ 46] = -18'sd    857;
assign PRECOMP_P1[ 47] = -18'sd    780;
assign PRECOMP_P1[ 48] = -18'sd    163;
assign PRECOMP_P1[ 49] =  18'sd    699;
assign PRECOMP_P1[ 50] =  18'sd   1290;
assign PRECOMP_P1[ 51] =  18'sd   1149;
assign PRECOMP_P1[ 52] =  18'sd    172;
assign PRECOMP_P1[ 53] = -18'sd   1232;
assign PRECOMP_P1[ 54] = -18'sd   2256;
assign PRECOMP_P1[ 55] = -18'sd   2055;
assign PRECOMP_P1[ 56] = -18'sd    177;
assign PRECOMP_P1[ 57] =  18'sd   3130;
assign PRECOMP_P1[ 58] =  18'sd   6933;
assign PRECOMP_P1[ 59] =  18'sd   9954;
assign PRECOMP_P1[ 60] =  18'sd  11103;
assign PRECOMP_P1[ 61] =  18'sd   9954;
assign PRECOMP_P1[ 62] =  18'sd   6933;
assign PRECOMP_P1[ 63] =  18'sd   3130;
assign PRECOMP_P1[ 64] = -18'sd    177;
assign PRECOMP_P1[ 65] = -18'sd   2055;
assign PRECOMP_P1[ 66] = -18'sd   2256;
assign PRECOMP_P1[ 67] = -18'sd   1232;
assign PRECOMP_P1[ 68] =  18'sd    172;
assign PRECOMP_P1[ 69] =  18'sd   1149;
assign PRECOMP_P1[ 70] =  18'sd   1290;
assign PRECOMP_P1[ 71] =  18'sd    699;
assign PRECOMP_P1[ 72] = -18'sd    163;
assign PRECOMP_P1[ 73] = -18'sd    780;
assign PRECOMP_P1[ 74] = -18'sd    857;
assign PRECOMP_P1[ 75] = -18'sd    443;
assign PRECOMP_P1[ 76] =  18'sd    152;
assign PRECOMP_P1[ 77] =  18'sd    570;
assign PRECOMP_P1[ 78] =  18'sd    604;
assign PRECOMP_P1[ 79] =  18'sd    292;
assign PRECOMP_P1[ 80] = -18'sd    139;
assign PRECOMP_P1[ 81] = -18'sd    429;
assign PRECOMP_P1[ 82] = -18'sd    436;
assign PRECOMP_P1[ 83] = -18'sd    194;
assign PRECOMP_P1[ 84] =  18'sd    123;
assign PRECOMP_P1[ 85] =  18'sd    327;
assign PRECOMP_P1[ 86] =  18'sd    316;
assign PRECOMP_P1[ 87] =  18'sd    127;
assign PRECOMP_P1[ 88] = -18'sd    107;
assign PRECOMP_P1[ 89] = -18'sd    248;
assign PRECOMP_P1[ 90] = -18'sd    228;
assign PRECOMP_P1[ 91] = -18'sd     81;
assign PRECOMP_P1[ 92] =  18'sd     91;
assign PRECOMP_P1[ 93] =  18'sd    186;
assign PRECOMP_P1[ 94] =  18'sd    161;
assign PRECOMP_P1[ 95] =  18'sd     49;
assign PRECOMP_P1[ 96] = -18'sd     75;
assign PRECOMP_P1[ 97] = -18'sd    137;
assign PRECOMP_P1[ 98] = -18'sd    112;
assign PRECOMP_P1[ 99] = -18'sd     27;
assign PRECOMP_P1[100] =  18'sd     60;
assign PRECOMP_P1[101] =  18'sd     99;
assign PRECOMP_P1[102] =  18'sd     75;
assign PRECOMP_P1[103] =  18'sd     12;
assign PRECOMP_P1[104] = -18'sd     46;
assign PRECOMP_P1[105] = -18'sd     69;
assign PRECOMP_P1[106] = -18'sd     48;
assign PRECOMP_P1[107] = -18'sd      4;
assign PRECOMP_P1[108] =  18'sd     34;
assign PRECOMP_P1[109] =  18'sd     46;
assign PRECOMP_P1[110] =  18'sd     29;
assign PRECOMP_P1[111] = -18'sd      1;
assign PRECOMP_P1[112] = -18'sd     24;
assign PRECOMP_P1[113] = -18'sd     29;
assign PRECOMP_P1[114] = -18'sd     16;
assign PRECOMP_P1[115] =  18'sd      3;
assign PRECOMP_P1[116] =  18'sd     16;
assign PRECOMP_P1[117] =  18'sd     17;
assign PRECOMP_P1[118] =  18'sd      8;
assign PRECOMP_P1[119] = -18'sd      3;
assign PRECOMP_P1[120] = -18'sd     10;



//TX Filter 18'sd N1 LUT Coefficients (headroom)
assign PRECOMP_N1[  0] =  18'sd     10;
assign PRECOMP_N1[  1] =  18'sd      3;
assign PRECOMP_N1[  2] = -18'sd      8;
assign PRECOMP_N1[  3] = -18'sd     17;
assign PRECOMP_N1[  4] = -18'sd     16;
assign PRECOMP_N1[  5] = -18'sd      3;
assign PRECOMP_N1[  6] =  18'sd     16;
assign PRECOMP_N1[  7] =  18'sd     29;
assign PRECOMP_N1[  8] =  18'sd     24;
assign PRECOMP_N1[  9] =  18'sd      1;
assign PRECOMP_N1[ 10] = -18'sd     29;
assign PRECOMP_N1[ 11] = -18'sd     46;
assign PRECOMP_N1[ 12] = -18'sd     34;
assign PRECOMP_N1[ 13] =  18'sd      4;
assign PRECOMP_N1[ 14] =  18'sd     48;
assign PRECOMP_N1[ 15] =  18'sd     69;
assign PRECOMP_N1[ 16] =  18'sd     46;
assign PRECOMP_N1[ 17] = -18'sd     12;
assign PRECOMP_N1[ 18] = -18'sd     75;
assign PRECOMP_N1[ 19] = -18'sd     99;
assign PRECOMP_N1[ 20] = -18'sd     60;
assign PRECOMP_N1[ 21] =  18'sd     27;
assign PRECOMP_N1[ 22] =  18'sd    112;
assign PRECOMP_N1[ 23] =  18'sd    137;
assign PRECOMP_N1[ 24] =  18'sd     75;
assign PRECOMP_N1[ 25] = -18'sd     49;
assign PRECOMP_N1[ 26] = -18'sd    161;
assign PRECOMP_N1[ 27] = -18'sd    186;
assign PRECOMP_N1[ 28] = -18'sd     91;
assign PRECOMP_N1[ 29] =  18'sd     81;
assign PRECOMP_N1[ 30] =  18'sd    228;
assign PRECOMP_N1[ 31] =  18'sd    248;
assign PRECOMP_N1[ 32] =  18'sd    107;
assign PRECOMP_N1[ 33] = -18'sd    127;
assign PRECOMP_N1[ 34] = -18'sd    316;
assign PRECOMP_N1[ 35] = -18'sd    327;
assign PRECOMP_N1[ 36] = -18'sd    123;
assign PRECOMP_N1[ 37] =  18'sd    194;
assign PRECOMP_N1[ 38] =  18'sd    436;
assign PRECOMP_N1[ 39] =  18'sd    429;
assign PRECOMP_N1[ 40] =  18'sd    139;
assign PRECOMP_N1[ 41] = -18'sd    292;
assign PRECOMP_N1[ 42] = -18'sd    604;
assign PRECOMP_N1[ 43] = -18'sd    570;
assign PRECOMP_N1[ 44] = -18'sd    152;
assign PRECOMP_N1[ 45] =  18'sd    443;
assign PRECOMP_N1[ 46] =  18'sd    857;
assign PRECOMP_N1[ 47] =  18'sd    780;
assign PRECOMP_N1[ 48] =  18'sd    163;
assign PRECOMP_N1[ 49] = -18'sd    699;
assign PRECOMP_N1[ 50] = -18'sd   1290;
assign PRECOMP_N1[ 51] = -18'sd   1149;
assign PRECOMP_N1[ 52] = -18'sd    172;
assign PRECOMP_N1[ 53] =  18'sd   1232;
assign PRECOMP_N1[ 54] =  18'sd   2256;
assign PRECOMP_N1[ 55] =  18'sd   2055;
assign PRECOMP_N1[ 56] =  18'sd    177;
assign PRECOMP_N1[ 57] = -18'sd   3130;
assign PRECOMP_N1[ 58] = -18'sd   6933;
assign PRECOMP_N1[ 59] = -18'sd   9954;
assign PRECOMP_N1[ 60] = -18'sd  11103;
assign PRECOMP_N1[ 61] = -18'sd   9954;
assign PRECOMP_N1[ 62] = -18'sd   6933;
assign PRECOMP_N1[ 63] = -18'sd   3130;
assign PRECOMP_N1[ 64] =  18'sd    177;
assign PRECOMP_N1[ 65] =  18'sd   2055;
assign PRECOMP_N1[ 66] =  18'sd   2256;
assign PRECOMP_N1[ 67] =  18'sd   1232;
assign PRECOMP_N1[ 68] = -18'sd    172;
assign PRECOMP_N1[ 69] = -18'sd   1149;
assign PRECOMP_N1[ 70] = -18'sd   1290;
assign PRECOMP_N1[ 71] = -18'sd    699;
assign PRECOMP_N1[ 72] =  18'sd    163;
assign PRECOMP_N1[ 73] =  18'sd    780;
assign PRECOMP_N1[ 74] =  18'sd    857;
assign PRECOMP_N1[ 75] =  18'sd    443;
assign PRECOMP_N1[ 76] = -18'sd    152;
assign PRECOMP_N1[ 77] = -18'sd    570;
assign PRECOMP_N1[ 78] = -18'sd    604;
assign PRECOMP_N1[ 79] = -18'sd    292;
assign PRECOMP_N1[ 80] =  18'sd    139;
assign PRECOMP_N1[ 81] =  18'sd    429;
assign PRECOMP_N1[ 82] =  18'sd    436;
assign PRECOMP_N1[ 83] =  18'sd    194;
assign PRECOMP_N1[ 84] = -18'sd    123;
assign PRECOMP_N1[ 85] = -18'sd    327;
assign PRECOMP_N1[ 86] = -18'sd    316;
assign PRECOMP_N1[ 87] = -18'sd    127;
assign PRECOMP_N1[ 88] =  18'sd    107;
assign PRECOMP_N1[ 89] =  18'sd    248;
assign PRECOMP_N1[ 90] =  18'sd    228;
assign PRECOMP_N1[ 91] =  18'sd     81;
assign PRECOMP_N1[ 92] = -18'sd     91;
assign PRECOMP_N1[ 93] = -18'sd    186;
assign PRECOMP_N1[ 94] = -18'sd    161;
assign PRECOMP_N1[ 95] = -18'sd     49;
assign PRECOMP_N1[ 96] =  18'sd     75;
assign PRECOMP_N1[ 97] =  18'sd    137;
assign PRECOMP_N1[ 98] =  18'sd    112;
assign PRECOMP_N1[ 99] =  18'sd     27;
assign PRECOMP_N1[100] = -18'sd     60;
assign PRECOMP_N1[101] = -18'sd     99;
assign PRECOMP_N1[102] = -18'sd     75;
assign PRECOMP_N1[103] = -18'sd     12;
assign PRECOMP_N1[104] =  18'sd     46;
assign PRECOMP_N1[105] =  18'sd     69;
assign PRECOMP_N1[106] =  18'sd     48;
assign PRECOMP_N1[107] =  18'sd      4;
assign PRECOMP_N1[108] = -18'sd     34;
assign PRECOMP_N1[109] = -18'sd     46;
assign PRECOMP_N1[110] = -18'sd     29;
assign PRECOMP_N1[111] =  18'sd      1;
assign PRECOMP_N1[112] =  18'sd     24;
assign PRECOMP_N1[113] =  18'sd     29;
assign PRECOMP_N1[114] =  18'sd     16;
assign PRECOMP_N1[115] = -18'sd      3;
assign PRECOMP_N1[116] = -18'sd     16;
assign PRECOMP_N1[117] = -18'sd     17;
assign PRECOMP_N1[118] = -18'sd      8;
assign PRECOMP_N1[119] =  18'sd      3;
assign PRECOMP_N1[120] =  18'sd     10;



//TX Filter 18'sd N2 LUT Coefficients (headroom)
assign PRECOMP_N2[  0] =  18'sd     29;
assign PRECOMP_N2[  1] =  18'sd     10;
assign PRECOMP_N2[  2] = -18'sd     24;
assign PRECOMP_N2[  3] = -18'sd     51;
assign PRECOMP_N2[  4] = -18'sd     48;
assign PRECOMP_N2[  5] = -18'sd      9;
assign PRECOMP_N2[  6] =  18'sd     49;
assign PRECOMP_N2[  7] =  18'sd     87;
assign PRECOMP_N2[  8] =  18'sd     73;
assign PRECOMP_N2[  9] =  18'sd      3;
assign PRECOMP_N2[ 10] = -18'sd     87;
assign PRECOMP_N2[ 11] = -18'sd    137;
assign PRECOMP_N2[ 12] = -18'sd    103;
assign PRECOMP_N2[ 13] =  18'sd     11;
assign PRECOMP_N2[ 14] =  18'sd    144;
assign PRECOMP_N2[ 15] =  18'sd    205;
assign PRECOMP_N2[ 16] =  18'sd    139;
assign PRECOMP_N2[ 17] = -18'sd     37;
assign PRECOMP_N2[ 18] = -18'sd    224;
assign PRECOMP_N2[ 19] = -18'sd    295;
assign PRECOMP_N2[ 20] = -18'sd    180;
assign PRECOMP_N2[ 21] =  18'sd     80;
assign PRECOMP_N2[ 22] =  18'sd    334;
assign PRECOMP_N2[ 23] =  18'sd    410;
assign PRECOMP_N2[ 24] =  18'sd    225;
assign PRECOMP_N2[ 25] = -18'sd    145;
assign PRECOMP_N2[ 26] = -18'sd    483;
assign PRECOMP_N2[ 27] = -18'sd    557;
assign PRECOMP_N2[ 28] = -18'sd    272;
assign PRECOMP_N2[ 29] =  18'sd    242;
assign PRECOMP_N2[ 30] =  18'sd    682;
assign PRECOMP_N2[ 31] =  18'sd    742;
assign PRECOMP_N2[ 32] =  18'sd    321;
assign PRECOMP_N2[ 33] = -18'sd    381;
assign PRECOMP_N2[ 34] = -18'sd    946;
assign PRECOMP_N2[ 35] = -18'sd    978;
assign PRECOMP_N2[ 36] = -18'sd    370;
assign PRECOMP_N2[ 37] =  18'sd    582;
assign PRECOMP_N2[ 38] =  18'sd   1305;
assign PRECOMP_N2[ 39] =  18'sd   1286;
assign PRECOMP_N2[ 40] =  18'sd    415;
assign PRECOMP_N2[ 41] = -18'sd    876;
assign PRECOMP_N2[ 42] = -18'sd   1808;
assign PRECOMP_N2[ 43] = -18'sd   1706;
assign PRECOMP_N2[ 44] = -18'sd    456;
assign PRECOMP_N2[ 45] =  18'sd   1327;
assign PRECOMP_N2[ 46] =  18'sd   2565;
assign PRECOMP_N2[ 47] =  18'sd   2335;
assign PRECOMP_N2[ 48] =  18'sd    490;
assign PRECOMP_N2[ 49] = -18'sd   2093;
assign PRECOMP_N2[ 50] = -18'sd   3863;
assign PRECOMP_N2[ 51] = -18'sd   3439;
assign PRECOMP_N2[ 52] = -18'sd    515;
assign PRECOMP_N2[ 53] =  18'sd   3687;
assign PRECOMP_N2[ 54] =  18'sd   6756;
assign PRECOMP_N2[ 55] =  18'sd   6153;
assign PRECOMP_N2[ 56] =  18'sd    531;
assign PRECOMP_N2[ 57] = -18'sd   9372;
assign PRECOMP_N2[ 58] = -18'sd  20759;
assign PRECOMP_N2[ 59] = -18'sd  29802;
assign PRECOMP_N2[ 60] = -18'sd  33241;
assign PRECOMP_N2[ 61] = -18'sd  29802;
assign PRECOMP_N2[ 62] = -18'sd  20759;
assign PRECOMP_N2[ 63] = -18'sd   9372;
assign PRECOMP_N2[ 64] =  18'sd    531;
assign PRECOMP_N2[ 65] =  18'sd   6153;
assign PRECOMP_N2[ 66] =  18'sd   6756;
assign PRECOMP_N2[ 67] =  18'sd   3687;
assign PRECOMP_N2[ 68] = -18'sd    515;
assign PRECOMP_N2[ 69] = -18'sd   3439;
assign PRECOMP_N2[ 70] = -18'sd   3863;
assign PRECOMP_N2[ 71] = -18'sd   2093;
assign PRECOMP_N2[ 72] =  18'sd    490;
assign PRECOMP_N2[ 73] =  18'sd   2335;
assign PRECOMP_N2[ 74] =  18'sd   2565;
assign PRECOMP_N2[ 75] =  18'sd   1327;
assign PRECOMP_N2[ 76] = -18'sd    456;
assign PRECOMP_N2[ 77] = -18'sd   1706;
assign PRECOMP_N2[ 78] = -18'sd   1808;
assign PRECOMP_N2[ 79] = -18'sd    876;
assign PRECOMP_N2[ 80] =  18'sd    415;
assign PRECOMP_N2[ 81] =  18'sd   1286;
assign PRECOMP_N2[ 82] =  18'sd   1305;
assign PRECOMP_N2[ 83] =  18'sd    582;
assign PRECOMP_N2[ 84] = -18'sd    370;
assign PRECOMP_N2[ 85] = -18'sd    978;
assign PRECOMP_N2[ 86] = -18'sd    946;
assign PRECOMP_N2[ 87] = -18'sd    381;
assign PRECOMP_N2[ 88] =  18'sd    321;
assign PRECOMP_N2[ 89] =  18'sd    742;
assign PRECOMP_N2[ 90] =  18'sd    682;
assign PRECOMP_N2[ 91] =  18'sd    242;
assign PRECOMP_N2[ 92] = -18'sd    272;
assign PRECOMP_N2[ 93] = -18'sd    557;
assign PRECOMP_N2[ 94] = -18'sd    483;
assign PRECOMP_N2[ 95] = -18'sd    145;
assign PRECOMP_N2[ 96] =  18'sd    225;
assign PRECOMP_N2[ 97] =  18'sd    410;
assign PRECOMP_N2[ 98] =  18'sd    334;
assign PRECOMP_N2[ 99] =  18'sd     80;
assign PRECOMP_N2[100] = -18'sd    180;
assign PRECOMP_N2[101] = -18'sd    295;
assign PRECOMP_N2[102] = -18'sd    224;
assign PRECOMP_N2[103] = -18'sd     37;
assign PRECOMP_N2[104] =  18'sd    139;
assign PRECOMP_N2[105] =  18'sd    205;
assign PRECOMP_N2[106] =  18'sd    144;
assign PRECOMP_N2[107] =  18'sd     11;
assign PRECOMP_N2[108] = -18'sd    103;
assign PRECOMP_N2[109] = -18'sd    137;
assign PRECOMP_N2[110] = -18'sd     87;
assign PRECOMP_N2[111] =  18'sd      3;
assign PRECOMP_N2[112] =  18'sd     73;
assign PRECOMP_N2[113] =  18'sd     87;
assign PRECOMP_N2[114] =  18'sd     49;
assign PRECOMP_N2[115] = -18'sd      9;
assign PRECOMP_N2[116] = -18'sd     48;
assign PRECOMP_N2[117] = -18'sd     51;
assign PRECOMP_N2[118] = -18'sd     24;
assign PRECOMP_N2[119] =  18'sd     10;
assign PRECOMP_N2[120] =  18'sd     29;

