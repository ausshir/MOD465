
//Halfband Filter 18'sd Multiplier Coefficients (headroom)
assign coef[  0] =  18'sd    391;
assign coef[  1] =  18'sd      0;
assign coef[  2] = -18'sd  10430;
assign coef[  3] =  18'sd      0;
assign coef[  4] =  18'sd  75478;
assign coef[  5] =  18'sd 131072;
