
//TX Filter 18'sd P2 LUT Coefficients (headroom)
assign PRECOMP_P2[  0] =  18'sd      3;
assign PRECOMP_P2[  1] = -18'sd      7;
assign PRECOMP_P2[  2] = -18'sd     12;
assign PRECOMP_P2[  3] = -18'sd      8;
assign PRECOMP_P2[  4] =  18'sd      2;
assign PRECOMP_P2[  5] =  18'sd     11;
assign PRECOMP_P2[  6] =  18'sd     12;
assign PRECOMP_P2[  7] =  18'sd      4;
assign PRECOMP_P2[  8] = -18'sd      7;
assign PRECOMP_P2[  9] = -18'sd     13;
assign PRECOMP_P2[ 10] = -18'sd     10;
assign PRECOMP_P2[ 11] =  18'sd      1;
assign PRECOMP_P2[ 12] =  18'sd     11;
assign PRECOMP_P2[ 13] =  18'sd     14;
assign PRECOMP_P2[ 14] =  18'sd      6;
assign PRECOMP_P2[ 15] = -18'sd      7;
assign PRECOMP_P2[ 16] = -18'sd     15;
assign PRECOMP_P2[ 17] = -18'sd     12;
assign PRECOMP_P2[ 18] =  18'sd      0;
assign PRECOMP_P2[ 19] =  18'sd     13;
assign PRECOMP_P2[ 20] =  18'sd     17;
assign PRECOMP_P2[ 21] =  18'sd      9;
assign PRECOMP_P2[ 22] = -18'sd      6;
assign PRECOMP_P2[ 23] = -18'sd     18;
assign PRECOMP_P2[ 24] = -18'sd     16;
assign PRECOMP_P2[ 25] = -18'sd      3;
assign PRECOMP_P2[ 26] =  18'sd     13;
assign PRECOMP_P2[ 27] =  18'sd     20;
assign PRECOMP_P2[ 28] =  18'sd     13;
assign PRECOMP_P2[ 29] = -18'sd      3;
assign PRECOMP_P2[ 30] = -18'sd     18;
assign PRECOMP_P2[ 31] = -18'sd     20;
assign PRECOMP_P2[ 32] = -18'sd      8;
assign PRECOMP_P2[ 33] =  18'sd     11;
assign PRECOMP_P2[ 34] =  18'sd     22;
assign PRECOMP_P2[ 35] =  18'sd     17;
assign PRECOMP_P2[ 36] =  18'sd      0;
assign PRECOMP_P2[ 37] = -18'sd     17;
assign PRECOMP_P2[ 38] = -18'sd     22;
assign PRECOMP_P2[ 39] = -18'sd     11;
assign PRECOMP_P2[ 40] =  18'sd      9;
assign PRECOMP_P2[ 41] =  18'sd     22;
assign PRECOMP_P2[ 42] =  18'sd     20;
assign PRECOMP_P2[ 43] =  18'sd      2;
assign PRECOMP_P2[ 44] = -18'sd     18;
assign PRECOMP_P2[ 45] = -18'sd     25;
assign PRECOMP_P2[ 46] = -18'sd     13;
assign PRECOMP_P2[ 47] =  18'sd      9;
assign PRECOMP_P2[ 48] =  18'sd     26;
assign PRECOMP_P2[ 49] =  18'sd     24;
assign PRECOMP_P2[ 50] =  18'sd      3;
assign PRECOMP_P2[ 51] = -18'sd     21;
assign PRECOMP_P2[ 52] = -18'sd     32;
assign PRECOMP_P2[ 53] = -18'sd     19;
assign PRECOMP_P2[ 54] =  18'sd      9;
assign PRECOMP_P2[ 55] =  18'sd     32;
assign PRECOMP_P2[ 56] =  18'sd     33;
assign PRECOMP_P2[ 57] =  18'sd     10;
assign PRECOMP_P2[ 58] = -18'sd     22;
assign PRECOMP_P2[ 59] = -18'sd     40;
assign PRECOMP_P2[ 60] = -18'sd     30;
assign PRECOMP_P2[ 61] =  18'sd      2;
assign PRECOMP_P2[ 62] =  18'sd     34;
assign PRECOMP_P2[ 63] =  18'sd     43;
assign PRECOMP_P2[ 64] =  18'sd     21;
assign PRECOMP_P2[ 65] = -18'sd     17;
assign PRECOMP_P2[ 66] = -18'sd     44;
assign PRECOMP_P2[ 67] = -18'sd     40;
assign PRECOMP_P2[ 68] = -18'sd      8;
assign PRECOMP_P2[ 69] =  18'sd     31;
assign PRECOMP_P2[ 70] =  18'sd     48;
assign PRECOMP_P2[ 71] =  18'sd     30;
assign PRECOMP_P2[ 72] = -18'sd     11;
assign PRECOMP_P2[ 73] = -18'sd     44;
assign PRECOMP_P2[ 74] = -18'sd     45;
assign PRECOMP_P2[ 75] = -18'sd     12;
assign PRECOMP_P2[ 76] =  18'sd     32;
assign PRECOMP_P2[ 77] =  18'sd     53;
assign PRECOMP_P2[ 78] =  18'sd     34;
assign PRECOMP_P2[ 79] = -18'sd     13;
assign PRECOMP_P2[ 80] = -18'sd     53;
assign PRECOMP_P2[ 81] = -18'sd     55;
assign PRECOMP_P2[ 82] = -18'sd     13;
assign PRECOMP_P2[ 83] =  18'sd     42;
assign PRECOMP_P2[ 84] =  18'sd     71;
assign PRECOMP_P2[ 85] =  18'sd     48;
assign PRECOMP_P2[ 86] = -18'sd     15;
assign PRECOMP_P2[ 87] = -18'sd     73;
assign PRECOMP_P2[ 88] = -18'sd     83;
assign PRECOMP_P2[ 89] = -18'sd     32;
assign PRECOMP_P2[ 90] =  18'sd     48;
assign PRECOMP_P2[ 91] =  18'sd    101;
assign PRECOMP_P2[ 92] =  18'sd     85;
assign PRECOMP_P2[ 93] =  18'sd      5;
assign PRECOMP_P2[ 94] = -18'sd     84;
assign PRECOMP_P2[ 95] = -18'sd    120;
assign PRECOMP_P2[ 96] = -18'sd     73;
assign PRECOMP_P2[ 97] =  18'sd     30;
assign PRECOMP_P2[ 98] =  18'sd    117;
assign PRECOMP_P2[ 99] =  18'sd    125;
assign PRECOMP_P2[100] =  18'sd     44;
assign PRECOMP_P2[101] = -18'sd     71;
assign PRECOMP_P2[102] = -18'sd    139;
assign PRECOMP_P2[103] = -18'sd    108;
assign PRECOMP_P2[104] =  18'sd      3;
assign PRECOMP_P2[105] =  18'sd    114;
assign PRECOMP_P2[106] =  18'sd    143;
assign PRECOMP_P2[107] =  18'sd     64;
assign PRECOMP_P2[108] = -18'sd     69;
assign PRECOMP_P2[109] = -18'sd    153;
assign PRECOMP_P2[110] = -18'sd    119;
assign PRECOMP_P2[111] =  18'sd     16;
assign PRECOMP_P2[112] =  18'sd    153;
assign PRECOMP_P2[113] =  18'sd    179;
assign PRECOMP_P2[114] =  18'sd     57;
assign PRECOMP_P2[115] = -18'sd    137;
assign PRECOMP_P2[116] = -18'sd    255;
assign PRECOMP_P2[117] = -18'sd    183;
assign PRECOMP_P2[118] =  18'sd     57;
assign PRECOMP_P2[119] =  18'sd    308;
assign PRECOMP_P2[120] =  18'sd    369;
assign PRECOMP_P2[121] =  18'sd    151;
assign PRECOMP_P2[122] = -18'sd    237;
assign PRECOMP_P2[123] = -18'sd    534;
assign PRECOMP_P2[124] = -18'sd    492;
assign PRECOMP_P2[125] = -18'sd     68;
assign PRECOMP_P2[126] =  18'sd    503;
assign PRECOMP_P2[127] =  18'sd    828;
assign PRECOMP_P2[128] =  18'sd    617;
assign PRECOMP_P2[129] = -18'sd     90;
assign PRECOMP_P2[130] = -18'sd    882;
assign PRECOMP_P2[131] = -18'sd   1208;
assign PRECOMP_P2[132] = -18'sd    738;
assign PRECOMP_P2[133] =  18'sd    357;
assign PRECOMP_P2[134] =  18'sd   1427;
assign PRECOMP_P2[135] =  18'sd   1713;
assign PRECOMP_P2[136] =  18'sd    848;
assign PRECOMP_P2[137] = -18'sd    801;
assign PRECOMP_P2[138] = -18'sd   2246;
assign PRECOMP_P2[139] = -18'sd   2432;
assign PRECOMP_P2[140] = -18'sd    942;
assign PRECOMP_P2[141] =  18'sd   1579;
assign PRECOMP_P2[142] =  18'sd   3622;
assign PRECOMP_P2[143] =  18'sd   3629;
assign PRECOMP_P2[144] =  18'sd   1013;
assign PRECOMP_P2[145] = -18'sd   3207;
assign PRECOMP_P2[146] = -18'sd   6607;
assign PRECOMP_P2[147] = -18'sd   6434;
assign PRECOMP_P2[148] = -18'sd   1057;
assign PRECOMP_P2[149] =  18'sd   8945;
assign PRECOMP_P2[150] =  18'sd  20712;
assign PRECOMP_P2[151] =  18'sd  30169;
assign PRECOMP_P2[152] =  18'sd  33785;
assign PRECOMP_P2[153] =  18'sd  30169;
assign PRECOMP_P2[154] =  18'sd  20712;
assign PRECOMP_P2[155] =  18'sd   8945;
assign PRECOMP_P2[156] = -18'sd   1057;
assign PRECOMP_P2[157] = -18'sd   6434;
assign PRECOMP_P2[158] = -18'sd   6607;
assign PRECOMP_P2[159] = -18'sd   3207;
assign PRECOMP_P2[160] =  18'sd   1013;
assign PRECOMP_P2[161] =  18'sd   3629;
assign PRECOMP_P2[162] =  18'sd   3622;
assign PRECOMP_P2[163] =  18'sd   1579;
assign PRECOMP_P2[164] = -18'sd    942;
assign PRECOMP_P2[165] = -18'sd   2432;
assign PRECOMP_P2[166] = -18'sd   2246;
assign PRECOMP_P2[167] = -18'sd    801;
assign PRECOMP_P2[168] =  18'sd    848;
assign PRECOMP_P2[169] =  18'sd   1713;
assign PRECOMP_P2[170] =  18'sd   1427;
assign PRECOMP_P2[171] =  18'sd    357;
assign PRECOMP_P2[172] = -18'sd    738;
assign PRECOMP_P2[173] = -18'sd   1208;
assign PRECOMP_P2[174] = -18'sd    882;
assign PRECOMP_P2[175] = -18'sd     90;
assign PRECOMP_P2[176] =  18'sd    617;
assign PRECOMP_P2[177] =  18'sd    828;
assign PRECOMP_P2[178] =  18'sd    503;
assign PRECOMP_P2[179] = -18'sd     68;
assign PRECOMP_P2[180] = -18'sd    492;
assign PRECOMP_P2[181] = -18'sd    534;
assign PRECOMP_P2[182] = -18'sd    237;
assign PRECOMP_P2[183] =  18'sd    151;
assign PRECOMP_P2[184] =  18'sd    369;
assign PRECOMP_P2[185] =  18'sd    308;
assign PRECOMP_P2[186] =  18'sd     57;
assign PRECOMP_P2[187] = -18'sd    183;
assign PRECOMP_P2[188] = -18'sd    255;
assign PRECOMP_P2[189] = -18'sd    137;
assign PRECOMP_P2[190] =  18'sd     57;
assign PRECOMP_P2[191] =  18'sd    179;
assign PRECOMP_P2[192] =  18'sd    153;
assign PRECOMP_P2[193] =  18'sd     16;
assign PRECOMP_P2[194] = -18'sd    119;
assign PRECOMP_P2[195] = -18'sd    153;
assign PRECOMP_P2[196] = -18'sd     69;
assign PRECOMP_P2[197] =  18'sd     64;
assign PRECOMP_P2[198] =  18'sd    143;
assign PRECOMP_P2[199] =  18'sd    114;
assign PRECOMP_P2[200] =  18'sd      3;
assign PRECOMP_P2[201] = -18'sd    108;
assign PRECOMP_P2[202] = -18'sd    139;
assign PRECOMP_P2[203] = -18'sd     71;
assign PRECOMP_P2[204] =  18'sd     44;
assign PRECOMP_P2[205] =  18'sd    125;
assign PRECOMP_P2[206] =  18'sd    117;
assign PRECOMP_P2[207] =  18'sd     30;
assign PRECOMP_P2[208] = -18'sd     73;
assign PRECOMP_P2[209] = -18'sd    120;
assign PRECOMP_P2[210] = -18'sd     84;
assign PRECOMP_P2[211] =  18'sd      5;
assign PRECOMP_P2[212] =  18'sd     85;
assign PRECOMP_P2[213] =  18'sd    101;
assign PRECOMP_P2[214] =  18'sd     48;
assign PRECOMP_P2[215] = -18'sd     32;
assign PRECOMP_P2[216] = -18'sd     83;
assign PRECOMP_P2[217] = -18'sd     73;
assign PRECOMP_P2[218] = -18'sd     15;
assign PRECOMP_P2[219] =  18'sd     48;
assign PRECOMP_P2[220] =  18'sd     71;
assign PRECOMP_P2[221] =  18'sd     42;
assign PRECOMP_P2[222] = -18'sd     13;
assign PRECOMP_P2[223] = -18'sd     55;
assign PRECOMP_P2[224] = -18'sd     53;
assign PRECOMP_P2[225] = -18'sd     13;
assign PRECOMP_P2[226] =  18'sd     34;
assign PRECOMP_P2[227] =  18'sd     53;
assign PRECOMP_P2[228] =  18'sd     32;
assign PRECOMP_P2[229] = -18'sd     12;
assign PRECOMP_P2[230] = -18'sd     45;
assign PRECOMP_P2[231] = -18'sd     44;
assign PRECOMP_P2[232] = -18'sd     11;
assign PRECOMP_P2[233] =  18'sd     30;
assign PRECOMP_P2[234] =  18'sd     48;
assign PRECOMP_P2[235] =  18'sd     31;
assign PRECOMP_P2[236] = -18'sd      8;
assign PRECOMP_P2[237] = -18'sd     40;
assign PRECOMP_P2[238] = -18'sd     44;
assign PRECOMP_P2[239] = -18'sd     17;
assign PRECOMP_P2[240] =  18'sd     21;
assign PRECOMP_P2[241] =  18'sd     43;
assign PRECOMP_P2[242] =  18'sd     34;
assign PRECOMP_P2[243] =  18'sd      2;
assign PRECOMP_P2[244] = -18'sd     30;
assign PRECOMP_P2[245] = -18'sd     40;
assign PRECOMP_P2[246] = -18'sd     22;
assign PRECOMP_P2[247] =  18'sd     10;
assign PRECOMP_P2[248] =  18'sd     33;
assign PRECOMP_P2[249] =  18'sd     32;
assign PRECOMP_P2[250] =  18'sd      9;
assign PRECOMP_P2[251] = -18'sd     19;
assign PRECOMP_P2[252] = -18'sd     32;
assign PRECOMP_P2[253] = -18'sd     21;
assign PRECOMP_P2[254] =  18'sd      3;
assign PRECOMP_P2[255] =  18'sd     24;
assign PRECOMP_P2[256] =  18'sd     26;
assign PRECOMP_P2[257] =  18'sd      9;
assign PRECOMP_P2[258] = -18'sd     13;
assign PRECOMP_P2[259] = -18'sd     25;
assign PRECOMP_P2[260] = -18'sd     18;
assign PRECOMP_P2[261] =  18'sd      2;
assign PRECOMP_P2[262] =  18'sd     20;
assign PRECOMP_P2[263] =  18'sd     22;
assign PRECOMP_P2[264] =  18'sd      9;
assign PRECOMP_P2[265] = -18'sd     11;
assign PRECOMP_P2[266] = -18'sd     22;
assign PRECOMP_P2[267] = -18'sd     17;
assign PRECOMP_P2[268] =  18'sd      0;
assign PRECOMP_P2[269] =  18'sd     17;
assign PRECOMP_P2[270] =  18'sd     22;
assign PRECOMP_P2[271] =  18'sd     11;
assign PRECOMP_P2[272] = -18'sd      8;
assign PRECOMP_P2[273] = -18'sd     20;
assign PRECOMP_P2[274] = -18'sd     18;
assign PRECOMP_P2[275] = -18'sd      3;
assign PRECOMP_P2[276] =  18'sd     13;
assign PRECOMP_P2[277] =  18'sd     20;
assign PRECOMP_P2[278] =  18'sd     13;
assign PRECOMP_P2[279] = -18'sd      3;
assign PRECOMP_P2[280] = -18'sd     16;
assign PRECOMP_P2[281] = -18'sd     18;
assign PRECOMP_P2[282] = -18'sd      6;
assign PRECOMP_P2[283] =  18'sd      9;
assign PRECOMP_P2[284] =  18'sd     17;
assign PRECOMP_P2[285] =  18'sd     13;
assign PRECOMP_P2[286] =  18'sd      0;
assign PRECOMP_P2[287] = -18'sd     12;
assign PRECOMP_P2[288] = -18'sd     15;
assign PRECOMP_P2[289] = -18'sd      7;
assign PRECOMP_P2[290] =  18'sd      6;
assign PRECOMP_P2[291] =  18'sd     14;
assign PRECOMP_P2[292] =  18'sd     11;
assign PRECOMP_P2[293] =  18'sd      1;
assign PRECOMP_P2[294] = -18'sd     10;
assign PRECOMP_P2[295] = -18'sd     13;
assign PRECOMP_P2[296] = -18'sd      7;
assign PRECOMP_P2[297] =  18'sd      4;
assign PRECOMP_P2[298] =  18'sd     12;
assign PRECOMP_P2[299] =  18'sd     11;
assign PRECOMP_P2[300] =  18'sd      2;
assign PRECOMP_P2[301] = -18'sd      8;
assign PRECOMP_P2[302] = -18'sd     12;
assign PRECOMP_P2[303] = -18'sd      7;
assign PRECOMP_P2[304] =  18'sd      3;



//TX Filter 18'sd P1 LUT Coefficients (headroom)
assign PRECOMP_P1[  0] =  18'sd      1;
assign PRECOMP_P1[  1] = -18'sd      2;
assign PRECOMP_P1[  2] = -18'sd      4;
assign PRECOMP_P1[  3] = -18'sd      3;
assign PRECOMP_P1[  4] =  18'sd      1;
assign PRECOMP_P1[  5] =  18'sd      4;
assign PRECOMP_P1[  6] =  18'sd      4;
assign PRECOMP_P1[  7] =  18'sd      1;
assign PRECOMP_P1[  8] = -18'sd      2;
assign PRECOMP_P1[  9] = -18'sd      4;
assign PRECOMP_P1[ 10] = -18'sd      3;
assign PRECOMP_P1[ 11] =  18'sd      0;
assign PRECOMP_P1[ 12] =  18'sd      4;
assign PRECOMP_P1[ 13] =  18'sd      5;
assign PRECOMP_P1[ 14] =  18'sd      2;
assign PRECOMP_P1[ 15] = -18'sd      2;
assign PRECOMP_P1[ 16] = -18'sd      5;
assign PRECOMP_P1[ 17] = -18'sd      4;
assign PRECOMP_P1[ 18] =  18'sd      0;
assign PRECOMP_P1[ 19] =  18'sd      4;
assign PRECOMP_P1[ 20] =  18'sd      6;
assign PRECOMP_P1[ 21] =  18'sd      3;
assign PRECOMP_P1[ 22] = -18'sd      2;
assign PRECOMP_P1[ 23] = -18'sd      6;
assign PRECOMP_P1[ 24] = -18'sd      5;
assign PRECOMP_P1[ 25] = -18'sd      1;
assign PRECOMP_P1[ 26] =  18'sd      4;
assign PRECOMP_P1[ 27] =  18'sd      7;
assign PRECOMP_P1[ 28] =  18'sd      4;
assign PRECOMP_P1[ 29] = -18'sd      1;
assign PRECOMP_P1[ 30] = -18'sd      6;
assign PRECOMP_P1[ 31] = -18'sd      7;
assign PRECOMP_P1[ 32] = -18'sd      3;
assign PRECOMP_P1[ 33] =  18'sd      4;
assign PRECOMP_P1[ 34] =  18'sd      7;
assign PRECOMP_P1[ 35] =  18'sd      6;
assign PRECOMP_P1[ 36] =  18'sd      0;
assign PRECOMP_P1[ 37] = -18'sd      6;
assign PRECOMP_P1[ 38] = -18'sd      7;
assign PRECOMP_P1[ 39] = -18'sd      4;
assign PRECOMP_P1[ 40] =  18'sd      3;
assign PRECOMP_P1[ 41] =  18'sd      7;
assign PRECOMP_P1[ 42] =  18'sd      7;
assign PRECOMP_P1[ 43] =  18'sd      1;
assign PRECOMP_P1[ 44] = -18'sd      6;
assign PRECOMP_P1[ 45] = -18'sd      8;
assign PRECOMP_P1[ 46] = -18'sd      4;
assign PRECOMP_P1[ 47] =  18'sd      3;
assign PRECOMP_P1[ 48] =  18'sd      9;
assign PRECOMP_P1[ 49] =  18'sd      8;
assign PRECOMP_P1[ 50] =  18'sd      1;
assign PRECOMP_P1[ 51] = -18'sd      7;
assign PRECOMP_P1[ 52] = -18'sd     11;
assign PRECOMP_P1[ 53] = -18'sd      6;
assign PRECOMP_P1[ 54] =  18'sd      3;
assign PRECOMP_P1[ 55] =  18'sd     11;
assign PRECOMP_P1[ 56] =  18'sd     11;
assign PRECOMP_P1[ 57] =  18'sd      3;
assign PRECOMP_P1[ 58] = -18'sd      7;
assign PRECOMP_P1[ 59] = -18'sd     13;
assign PRECOMP_P1[ 60] = -18'sd     10;
assign PRECOMP_P1[ 61] =  18'sd      1;
assign PRECOMP_P1[ 62] =  18'sd     12;
assign PRECOMP_P1[ 63] =  18'sd     14;
assign PRECOMP_P1[ 64] =  18'sd      7;
assign PRECOMP_P1[ 65] = -18'sd      6;
assign PRECOMP_P1[ 66] = -18'sd     15;
assign PRECOMP_P1[ 67] = -18'sd     13;
assign PRECOMP_P1[ 68] = -18'sd      3;
assign PRECOMP_P1[ 69] =  18'sd     10;
assign PRECOMP_P1[ 70] =  18'sd     16;
assign PRECOMP_P1[ 71] =  18'sd     10;
assign PRECOMP_P1[ 72] = -18'sd      4;
assign PRECOMP_P1[ 73] = -18'sd     15;
assign PRECOMP_P1[ 74] = -18'sd     15;
assign PRECOMP_P1[ 75] = -18'sd      4;
assign PRECOMP_P1[ 76] =  18'sd     11;
assign PRECOMP_P1[ 77] =  18'sd     18;
assign PRECOMP_P1[ 78] =  18'sd     11;
assign PRECOMP_P1[ 79] = -18'sd      4;
assign PRECOMP_P1[ 80] = -18'sd     18;
assign PRECOMP_P1[ 81] = -18'sd     18;
assign PRECOMP_P1[ 82] = -18'sd      4;
assign PRECOMP_P1[ 83] =  18'sd     14;
assign PRECOMP_P1[ 84] =  18'sd     24;
assign PRECOMP_P1[ 85] =  18'sd     16;
assign PRECOMP_P1[ 86] = -18'sd      5;
assign PRECOMP_P1[ 87] = -18'sd     24;
assign PRECOMP_P1[ 88] = -18'sd     28;
assign PRECOMP_P1[ 89] = -18'sd     11;
assign PRECOMP_P1[ 90] =  18'sd     16;
assign PRECOMP_P1[ 91] =  18'sd     34;
assign PRECOMP_P1[ 92] =  18'sd     28;
assign PRECOMP_P1[ 93] =  18'sd      2;
assign PRECOMP_P1[ 94] = -18'sd     28;
assign PRECOMP_P1[ 95] = -18'sd     40;
assign PRECOMP_P1[ 96] = -18'sd     24;
assign PRECOMP_P1[ 97] =  18'sd     10;
assign PRECOMP_P1[ 98] =  18'sd     39;
assign PRECOMP_P1[ 99] =  18'sd     42;
assign PRECOMP_P1[100] =  18'sd     15;
assign PRECOMP_P1[101] = -18'sd     24;
assign PRECOMP_P1[102] = -18'sd     47;
assign PRECOMP_P1[103] = -18'sd     36;
assign PRECOMP_P1[104] =  18'sd      1;
assign PRECOMP_P1[105] =  18'sd     38;
assign PRECOMP_P1[106] =  18'sd     48;
assign PRECOMP_P1[107] =  18'sd     21;
assign PRECOMP_P1[108] = -18'sd     23;
assign PRECOMP_P1[109] = -18'sd     51;
assign PRECOMP_P1[110] = -18'sd     40;
assign PRECOMP_P1[111] =  18'sd      5;
assign PRECOMP_P1[112] =  18'sd     51;
assign PRECOMP_P1[113] =  18'sd     60;
assign PRECOMP_P1[114] =  18'sd     19;
assign PRECOMP_P1[115] = -18'sd     46;
assign PRECOMP_P1[116] = -18'sd     85;
assign PRECOMP_P1[117] = -18'sd     61;
assign PRECOMP_P1[118] =  18'sd     19;
assign PRECOMP_P1[119] =  18'sd    103;
assign PRECOMP_P1[120] =  18'sd    123;
assign PRECOMP_P1[121] =  18'sd     50;
assign PRECOMP_P1[122] = -18'sd     79;
assign PRECOMP_P1[123] = -18'sd    178;
assign PRECOMP_P1[124] = -18'sd    164;
assign PRECOMP_P1[125] = -18'sd     23;
assign PRECOMP_P1[126] =  18'sd    168;
assign PRECOMP_P1[127] =  18'sd    277;
assign PRECOMP_P1[128] =  18'sd    206;
assign PRECOMP_P1[129] = -18'sd     30;
assign PRECOMP_P1[130] = -18'sd    295;
assign PRECOMP_P1[131] = -18'sd    403;
assign PRECOMP_P1[132] = -18'sd    246;
assign PRECOMP_P1[133] =  18'sd    119;
assign PRECOMP_P1[134] =  18'sd    477;
assign PRECOMP_P1[135] =  18'sd    572;
assign PRECOMP_P1[136] =  18'sd    283;
assign PRECOMP_P1[137] = -18'sd    267;
assign PRECOMP_P1[138] = -18'sd    750;
assign PRECOMP_P1[139] = -18'sd    812;
assign PRECOMP_P1[140] = -18'sd    315;
assign PRECOMP_P1[141] =  18'sd    527;
assign PRECOMP_P1[142] =  18'sd   1210;
assign PRECOMP_P1[143] =  18'sd   1212;
assign PRECOMP_P1[144] =  18'sd    338;
assign PRECOMP_P1[145] = -18'sd   1071;
assign PRECOMP_P1[146] = -18'sd   2207;
assign PRECOMP_P1[147] = -18'sd   2149;
assign PRECOMP_P1[148] = -18'sd    353;
assign PRECOMP_P1[149] =  18'sd   2988;
assign PRECOMP_P1[150] =  18'sd   6918;
assign PRECOMP_P1[151] =  18'sd  10076;
assign PRECOMP_P1[152] =  18'sd  11284;
assign PRECOMP_P1[153] =  18'sd  10076;
assign PRECOMP_P1[154] =  18'sd   6918;
assign PRECOMP_P1[155] =  18'sd   2988;
assign PRECOMP_P1[156] = -18'sd    353;
assign PRECOMP_P1[157] = -18'sd   2149;
assign PRECOMP_P1[158] = -18'sd   2207;
assign PRECOMP_P1[159] = -18'sd   1071;
assign PRECOMP_P1[160] =  18'sd    338;
assign PRECOMP_P1[161] =  18'sd   1212;
assign PRECOMP_P1[162] =  18'sd   1210;
assign PRECOMP_P1[163] =  18'sd    527;
assign PRECOMP_P1[164] = -18'sd    315;
assign PRECOMP_P1[165] = -18'sd    812;
assign PRECOMP_P1[166] = -18'sd    750;
assign PRECOMP_P1[167] = -18'sd    267;
assign PRECOMP_P1[168] =  18'sd    283;
assign PRECOMP_P1[169] =  18'sd    572;
assign PRECOMP_P1[170] =  18'sd    477;
assign PRECOMP_P1[171] =  18'sd    119;
assign PRECOMP_P1[172] = -18'sd    246;
assign PRECOMP_P1[173] = -18'sd    403;
assign PRECOMP_P1[174] = -18'sd    295;
assign PRECOMP_P1[175] = -18'sd     30;
assign PRECOMP_P1[176] =  18'sd    206;
assign PRECOMP_P1[177] =  18'sd    277;
assign PRECOMP_P1[178] =  18'sd    168;
assign PRECOMP_P1[179] = -18'sd     23;
assign PRECOMP_P1[180] = -18'sd    164;
assign PRECOMP_P1[181] = -18'sd    178;
assign PRECOMP_P1[182] = -18'sd     79;
assign PRECOMP_P1[183] =  18'sd     50;
assign PRECOMP_P1[184] =  18'sd    123;
assign PRECOMP_P1[185] =  18'sd    103;
assign PRECOMP_P1[186] =  18'sd     19;
assign PRECOMP_P1[187] = -18'sd     61;
assign PRECOMP_P1[188] = -18'sd     85;
assign PRECOMP_P1[189] = -18'sd     46;
assign PRECOMP_P1[190] =  18'sd     19;
assign PRECOMP_P1[191] =  18'sd     60;
assign PRECOMP_P1[192] =  18'sd     51;
assign PRECOMP_P1[193] =  18'sd      5;
assign PRECOMP_P1[194] = -18'sd     40;
assign PRECOMP_P1[195] = -18'sd     51;
assign PRECOMP_P1[196] = -18'sd     23;
assign PRECOMP_P1[197] =  18'sd     21;
assign PRECOMP_P1[198] =  18'sd     48;
assign PRECOMP_P1[199] =  18'sd     38;
assign PRECOMP_P1[200] =  18'sd      1;
assign PRECOMP_P1[201] = -18'sd     36;
assign PRECOMP_P1[202] = -18'sd     47;
assign PRECOMP_P1[203] = -18'sd     24;
assign PRECOMP_P1[204] =  18'sd     15;
assign PRECOMP_P1[205] =  18'sd     42;
assign PRECOMP_P1[206] =  18'sd     39;
assign PRECOMP_P1[207] =  18'sd     10;
assign PRECOMP_P1[208] = -18'sd     24;
assign PRECOMP_P1[209] = -18'sd     40;
assign PRECOMP_P1[210] = -18'sd     28;
assign PRECOMP_P1[211] =  18'sd      2;
assign PRECOMP_P1[212] =  18'sd     28;
assign PRECOMP_P1[213] =  18'sd     34;
assign PRECOMP_P1[214] =  18'sd     16;
assign PRECOMP_P1[215] = -18'sd     11;
assign PRECOMP_P1[216] = -18'sd     28;
assign PRECOMP_P1[217] = -18'sd     24;
assign PRECOMP_P1[218] = -18'sd      5;
assign PRECOMP_P1[219] =  18'sd     16;
assign PRECOMP_P1[220] =  18'sd     24;
assign PRECOMP_P1[221] =  18'sd     14;
assign PRECOMP_P1[222] = -18'sd      4;
assign PRECOMP_P1[223] = -18'sd     18;
assign PRECOMP_P1[224] = -18'sd     18;
assign PRECOMP_P1[225] = -18'sd      4;
assign PRECOMP_P1[226] =  18'sd     11;
assign PRECOMP_P1[227] =  18'sd     18;
assign PRECOMP_P1[228] =  18'sd     11;
assign PRECOMP_P1[229] = -18'sd      4;
assign PRECOMP_P1[230] = -18'sd     15;
assign PRECOMP_P1[231] = -18'sd     15;
assign PRECOMP_P1[232] = -18'sd      4;
assign PRECOMP_P1[233] =  18'sd     10;
assign PRECOMP_P1[234] =  18'sd     16;
assign PRECOMP_P1[235] =  18'sd     10;
assign PRECOMP_P1[236] = -18'sd      3;
assign PRECOMP_P1[237] = -18'sd     13;
assign PRECOMP_P1[238] = -18'sd     15;
assign PRECOMP_P1[239] = -18'sd      6;
assign PRECOMP_P1[240] =  18'sd      7;
assign PRECOMP_P1[241] =  18'sd     14;
assign PRECOMP_P1[242] =  18'sd     12;
assign PRECOMP_P1[243] =  18'sd      1;
assign PRECOMP_P1[244] = -18'sd     10;
assign PRECOMP_P1[245] = -18'sd     13;
assign PRECOMP_P1[246] = -18'sd      7;
assign PRECOMP_P1[247] =  18'sd      3;
assign PRECOMP_P1[248] =  18'sd     11;
assign PRECOMP_P1[249] =  18'sd     11;
assign PRECOMP_P1[250] =  18'sd      3;
assign PRECOMP_P1[251] = -18'sd      6;
assign PRECOMP_P1[252] = -18'sd     11;
assign PRECOMP_P1[253] = -18'sd      7;
assign PRECOMP_P1[254] =  18'sd      1;
assign PRECOMP_P1[255] =  18'sd      8;
assign PRECOMP_P1[256] =  18'sd      9;
assign PRECOMP_P1[257] =  18'sd      3;
assign PRECOMP_P1[258] = -18'sd      4;
assign PRECOMP_P1[259] = -18'sd      8;
assign PRECOMP_P1[260] = -18'sd      6;
assign PRECOMP_P1[261] =  18'sd      1;
assign PRECOMP_P1[262] =  18'sd      7;
assign PRECOMP_P1[263] =  18'sd      7;
assign PRECOMP_P1[264] =  18'sd      3;
assign PRECOMP_P1[265] = -18'sd      4;
assign PRECOMP_P1[266] = -18'sd      7;
assign PRECOMP_P1[267] = -18'sd      6;
assign PRECOMP_P1[268] =  18'sd      0;
assign PRECOMP_P1[269] =  18'sd      6;
assign PRECOMP_P1[270] =  18'sd      7;
assign PRECOMP_P1[271] =  18'sd      4;
assign PRECOMP_P1[272] = -18'sd      3;
assign PRECOMP_P1[273] = -18'sd      7;
assign PRECOMP_P1[274] = -18'sd      6;
assign PRECOMP_P1[275] = -18'sd      1;
assign PRECOMP_P1[276] =  18'sd      4;
assign PRECOMP_P1[277] =  18'sd      7;
assign PRECOMP_P1[278] =  18'sd      4;
assign PRECOMP_P1[279] = -18'sd      1;
assign PRECOMP_P1[280] = -18'sd      5;
assign PRECOMP_P1[281] = -18'sd      6;
assign PRECOMP_P1[282] = -18'sd      2;
assign PRECOMP_P1[283] =  18'sd      3;
assign PRECOMP_P1[284] =  18'sd      6;
assign PRECOMP_P1[285] =  18'sd      4;
assign PRECOMP_P1[286] =  18'sd      0;
assign PRECOMP_P1[287] = -18'sd      4;
assign PRECOMP_P1[288] = -18'sd      5;
assign PRECOMP_P1[289] = -18'sd      2;
assign PRECOMP_P1[290] =  18'sd      2;
assign PRECOMP_P1[291] =  18'sd      5;
assign PRECOMP_P1[292] =  18'sd      4;
assign PRECOMP_P1[293] =  18'sd      0;
assign PRECOMP_P1[294] = -18'sd      3;
assign PRECOMP_P1[295] = -18'sd      4;
assign PRECOMP_P1[296] = -18'sd      2;
assign PRECOMP_P1[297] =  18'sd      1;
assign PRECOMP_P1[298] =  18'sd      4;
assign PRECOMP_P1[299] =  18'sd      4;
assign PRECOMP_P1[300] =  18'sd      1;
assign PRECOMP_P1[301] = -18'sd      3;
assign PRECOMP_P1[302] = -18'sd      4;
assign PRECOMP_P1[303] = -18'sd      2;
assign PRECOMP_P1[304] =  18'sd      1;



//TX Filter 18'sd N1 LUT Coefficients (headroom)
assign PRECOMP_N1[  0] = -18'sd      1;
assign PRECOMP_N1[  1] =  18'sd      2;
assign PRECOMP_N1[  2] =  18'sd      4;
assign PRECOMP_N1[  3] =  18'sd      3;
assign PRECOMP_N1[  4] = -18'sd      1;
assign PRECOMP_N1[  5] = -18'sd      4;
assign PRECOMP_N1[  6] = -18'sd      4;
assign PRECOMP_N1[  7] = -18'sd      1;
assign PRECOMP_N1[  8] =  18'sd      2;
assign PRECOMP_N1[  9] =  18'sd      4;
assign PRECOMP_N1[ 10] =  18'sd      3;
assign PRECOMP_N1[ 11] =  18'sd      0;
assign PRECOMP_N1[ 12] = -18'sd      4;
assign PRECOMP_N1[ 13] = -18'sd      5;
assign PRECOMP_N1[ 14] = -18'sd      2;
assign PRECOMP_N1[ 15] =  18'sd      2;
assign PRECOMP_N1[ 16] =  18'sd      5;
assign PRECOMP_N1[ 17] =  18'sd      4;
assign PRECOMP_N1[ 18] =  18'sd      0;
assign PRECOMP_N1[ 19] = -18'sd      4;
assign PRECOMP_N1[ 20] = -18'sd      6;
assign PRECOMP_N1[ 21] = -18'sd      3;
assign PRECOMP_N1[ 22] =  18'sd      2;
assign PRECOMP_N1[ 23] =  18'sd      6;
assign PRECOMP_N1[ 24] =  18'sd      5;
assign PRECOMP_N1[ 25] =  18'sd      1;
assign PRECOMP_N1[ 26] = -18'sd      4;
assign PRECOMP_N1[ 27] = -18'sd      7;
assign PRECOMP_N1[ 28] = -18'sd      4;
assign PRECOMP_N1[ 29] =  18'sd      1;
assign PRECOMP_N1[ 30] =  18'sd      6;
assign PRECOMP_N1[ 31] =  18'sd      7;
assign PRECOMP_N1[ 32] =  18'sd      3;
assign PRECOMP_N1[ 33] = -18'sd      4;
assign PRECOMP_N1[ 34] = -18'sd      7;
assign PRECOMP_N1[ 35] = -18'sd      6;
assign PRECOMP_N1[ 36] =  18'sd      0;
assign PRECOMP_N1[ 37] =  18'sd      6;
assign PRECOMP_N1[ 38] =  18'sd      7;
assign PRECOMP_N1[ 39] =  18'sd      4;
assign PRECOMP_N1[ 40] = -18'sd      3;
assign PRECOMP_N1[ 41] = -18'sd      7;
assign PRECOMP_N1[ 42] = -18'sd      7;
assign PRECOMP_N1[ 43] = -18'sd      1;
assign PRECOMP_N1[ 44] =  18'sd      6;
assign PRECOMP_N1[ 45] =  18'sd      8;
assign PRECOMP_N1[ 46] =  18'sd      4;
assign PRECOMP_N1[ 47] = -18'sd      3;
assign PRECOMP_N1[ 48] = -18'sd      9;
assign PRECOMP_N1[ 49] = -18'sd      8;
assign PRECOMP_N1[ 50] = -18'sd      1;
assign PRECOMP_N1[ 51] =  18'sd      7;
assign PRECOMP_N1[ 52] =  18'sd     11;
assign PRECOMP_N1[ 53] =  18'sd      6;
assign PRECOMP_N1[ 54] = -18'sd      3;
assign PRECOMP_N1[ 55] = -18'sd     11;
assign PRECOMP_N1[ 56] = -18'sd     11;
assign PRECOMP_N1[ 57] = -18'sd      3;
assign PRECOMP_N1[ 58] =  18'sd      7;
assign PRECOMP_N1[ 59] =  18'sd     13;
assign PRECOMP_N1[ 60] =  18'sd     10;
assign PRECOMP_N1[ 61] = -18'sd      1;
assign PRECOMP_N1[ 62] = -18'sd     12;
assign PRECOMP_N1[ 63] = -18'sd     14;
assign PRECOMP_N1[ 64] = -18'sd      7;
assign PRECOMP_N1[ 65] =  18'sd      6;
assign PRECOMP_N1[ 66] =  18'sd     15;
assign PRECOMP_N1[ 67] =  18'sd     13;
assign PRECOMP_N1[ 68] =  18'sd      3;
assign PRECOMP_N1[ 69] = -18'sd     10;
assign PRECOMP_N1[ 70] = -18'sd     16;
assign PRECOMP_N1[ 71] = -18'sd     10;
assign PRECOMP_N1[ 72] =  18'sd      4;
assign PRECOMP_N1[ 73] =  18'sd     15;
assign PRECOMP_N1[ 74] =  18'sd     15;
assign PRECOMP_N1[ 75] =  18'sd      4;
assign PRECOMP_N1[ 76] = -18'sd     11;
assign PRECOMP_N1[ 77] = -18'sd     18;
assign PRECOMP_N1[ 78] = -18'sd     11;
assign PRECOMP_N1[ 79] =  18'sd      4;
assign PRECOMP_N1[ 80] =  18'sd     18;
assign PRECOMP_N1[ 81] =  18'sd     18;
assign PRECOMP_N1[ 82] =  18'sd      4;
assign PRECOMP_N1[ 83] = -18'sd     14;
assign PRECOMP_N1[ 84] = -18'sd     24;
assign PRECOMP_N1[ 85] = -18'sd     16;
assign PRECOMP_N1[ 86] =  18'sd      5;
assign PRECOMP_N1[ 87] =  18'sd     24;
assign PRECOMP_N1[ 88] =  18'sd     28;
assign PRECOMP_N1[ 89] =  18'sd     11;
assign PRECOMP_N1[ 90] = -18'sd     16;
assign PRECOMP_N1[ 91] = -18'sd     34;
assign PRECOMP_N1[ 92] = -18'sd     28;
assign PRECOMP_N1[ 93] = -18'sd      2;
assign PRECOMP_N1[ 94] =  18'sd     28;
assign PRECOMP_N1[ 95] =  18'sd     40;
assign PRECOMP_N1[ 96] =  18'sd     24;
assign PRECOMP_N1[ 97] = -18'sd     10;
assign PRECOMP_N1[ 98] = -18'sd     39;
assign PRECOMP_N1[ 99] = -18'sd     42;
assign PRECOMP_N1[100] = -18'sd     15;
assign PRECOMP_N1[101] =  18'sd     24;
assign PRECOMP_N1[102] =  18'sd     47;
assign PRECOMP_N1[103] =  18'sd     36;
assign PRECOMP_N1[104] = -18'sd      1;
assign PRECOMP_N1[105] = -18'sd     38;
assign PRECOMP_N1[106] = -18'sd     48;
assign PRECOMP_N1[107] = -18'sd     21;
assign PRECOMP_N1[108] =  18'sd     23;
assign PRECOMP_N1[109] =  18'sd     51;
assign PRECOMP_N1[110] =  18'sd     40;
assign PRECOMP_N1[111] = -18'sd      5;
assign PRECOMP_N1[112] = -18'sd     51;
assign PRECOMP_N1[113] = -18'sd     60;
assign PRECOMP_N1[114] = -18'sd     19;
assign PRECOMP_N1[115] =  18'sd     46;
assign PRECOMP_N1[116] =  18'sd     85;
assign PRECOMP_N1[117] =  18'sd     61;
assign PRECOMP_N1[118] = -18'sd     19;
assign PRECOMP_N1[119] = -18'sd    103;
assign PRECOMP_N1[120] = -18'sd    123;
assign PRECOMP_N1[121] = -18'sd     50;
assign PRECOMP_N1[122] =  18'sd     79;
assign PRECOMP_N1[123] =  18'sd    178;
assign PRECOMP_N1[124] =  18'sd    164;
assign PRECOMP_N1[125] =  18'sd     23;
assign PRECOMP_N1[126] = -18'sd    168;
assign PRECOMP_N1[127] = -18'sd    277;
assign PRECOMP_N1[128] = -18'sd    206;
assign PRECOMP_N1[129] =  18'sd     30;
assign PRECOMP_N1[130] =  18'sd    295;
assign PRECOMP_N1[131] =  18'sd    403;
assign PRECOMP_N1[132] =  18'sd    246;
assign PRECOMP_N1[133] = -18'sd    119;
assign PRECOMP_N1[134] = -18'sd    477;
assign PRECOMP_N1[135] = -18'sd    572;
assign PRECOMP_N1[136] = -18'sd    283;
assign PRECOMP_N1[137] =  18'sd    267;
assign PRECOMP_N1[138] =  18'sd    750;
assign PRECOMP_N1[139] =  18'sd    812;
assign PRECOMP_N1[140] =  18'sd    315;
assign PRECOMP_N1[141] = -18'sd    527;
assign PRECOMP_N1[142] = -18'sd   1210;
assign PRECOMP_N1[143] = -18'sd   1212;
assign PRECOMP_N1[144] = -18'sd    338;
assign PRECOMP_N1[145] =  18'sd   1071;
assign PRECOMP_N1[146] =  18'sd   2207;
assign PRECOMP_N1[147] =  18'sd   2149;
assign PRECOMP_N1[148] =  18'sd    353;
assign PRECOMP_N1[149] = -18'sd   2988;
assign PRECOMP_N1[150] = -18'sd   6918;
assign PRECOMP_N1[151] = -18'sd  10076;
assign PRECOMP_N1[152] = -18'sd  11284;
assign PRECOMP_N1[153] = -18'sd  10076;
assign PRECOMP_N1[154] = -18'sd   6918;
assign PRECOMP_N1[155] = -18'sd   2988;
assign PRECOMP_N1[156] =  18'sd    353;
assign PRECOMP_N1[157] =  18'sd   2149;
assign PRECOMP_N1[158] =  18'sd   2207;
assign PRECOMP_N1[159] =  18'sd   1071;
assign PRECOMP_N1[160] = -18'sd    338;
assign PRECOMP_N1[161] = -18'sd   1212;
assign PRECOMP_N1[162] = -18'sd   1210;
assign PRECOMP_N1[163] = -18'sd    527;
assign PRECOMP_N1[164] =  18'sd    315;
assign PRECOMP_N1[165] =  18'sd    812;
assign PRECOMP_N1[166] =  18'sd    750;
assign PRECOMP_N1[167] =  18'sd    267;
assign PRECOMP_N1[168] = -18'sd    283;
assign PRECOMP_N1[169] = -18'sd    572;
assign PRECOMP_N1[170] = -18'sd    477;
assign PRECOMP_N1[171] = -18'sd    119;
assign PRECOMP_N1[172] =  18'sd    246;
assign PRECOMP_N1[173] =  18'sd    403;
assign PRECOMP_N1[174] =  18'sd    295;
assign PRECOMP_N1[175] =  18'sd     30;
assign PRECOMP_N1[176] = -18'sd    206;
assign PRECOMP_N1[177] = -18'sd    277;
assign PRECOMP_N1[178] = -18'sd    168;
assign PRECOMP_N1[179] =  18'sd     23;
assign PRECOMP_N1[180] =  18'sd    164;
assign PRECOMP_N1[181] =  18'sd    178;
assign PRECOMP_N1[182] =  18'sd     79;
assign PRECOMP_N1[183] = -18'sd     50;
assign PRECOMP_N1[184] = -18'sd    123;
assign PRECOMP_N1[185] = -18'sd    103;
assign PRECOMP_N1[186] = -18'sd     19;
assign PRECOMP_N1[187] =  18'sd     61;
assign PRECOMP_N1[188] =  18'sd     85;
assign PRECOMP_N1[189] =  18'sd     46;
assign PRECOMP_N1[190] = -18'sd     19;
assign PRECOMP_N1[191] = -18'sd     60;
assign PRECOMP_N1[192] = -18'sd     51;
assign PRECOMP_N1[193] = -18'sd      5;
assign PRECOMP_N1[194] =  18'sd     40;
assign PRECOMP_N1[195] =  18'sd     51;
assign PRECOMP_N1[196] =  18'sd     23;
assign PRECOMP_N1[197] = -18'sd     21;
assign PRECOMP_N1[198] = -18'sd     48;
assign PRECOMP_N1[199] = -18'sd     38;
assign PRECOMP_N1[200] = -18'sd      1;
assign PRECOMP_N1[201] =  18'sd     36;
assign PRECOMP_N1[202] =  18'sd     47;
assign PRECOMP_N1[203] =  18'sd     24;
assign PRECOMP_N1[204] = -18'sd     15;
assign PRECOMP_N1[205] = -18'sd     42;
assign PRECOMP_N1[206] = -18'sd     39;
assign PRECOMP_N1[207] = -18'sd     10;
assign PRECOMP_N1[208] =  18'sd     24;
assign PRECOMP_N1[209] =  18'sd     40;
assign PRECOMP_N1[210] =  18'sd     28;
assign PRECOMP_N1[211] = -18'sd      2;
assign PRECOMP_N1[212] = -18'sd     28;
assign PRECOMP_N1[213] = -18'sd     34;
assign PRECOMP_N1[214] = -18'sd     16;
assign PRECOMP_N1[215] =  18'sd     11;
assign PRECOMP_N1[216] =  18'sd     28;
assign PRECOMP_N1[217] =  18'sd     24;
assign PRECOMP_N1[218] =  18'sd      5;
assign PRECOMP_N1[219] = -18'sd     16;
assign PRECOMP_N1[220] = -18'sd     24;
assign PRECOMP_N1[221] = -18'sd     14;
assign PRECOMP_N1[222] =  18'sd      4;
assign PRECOMP_N1[223] =  18'sd     18;
assign PRECOMP_N1[224] =  18'sd     18;
assign PRECOMP_N1[225] =  18'sd      4;
assign PRECOMP_N1[226] = -18'sd     11;
assign PRECOMP_N1[227] = -18'sd     18;
assign PRECOMP_N1[228] = -18'sd     11;
assign PRECOMP_N1[229] =  18'sd      4;
assign PRECOMP_N1[230] =  18'sd     15;
assign PRECOMP_N1[231] =  18'sd     15;
assign PRECOMP_N1[232] =  18'sd      4;
assign PRECOMP_N1[233] = -18'sd     10;
assign PRECOMP_N1[234] = -18'sd     16;
assign PRECOMP_N1[235] = -18'sd     10;
assign PRECOMP_N1[236] =  18'sd      3;
assign PRECOMP_N1[237] =  18'sd     13;
assign PRECOMP_N1[238] =  18'sd     15;
assign PRECOMP_N1[239] =  18'sd      6;
assign PRECOMP_N1[240] = -18'sd      7;
assign PRECOMP_N1[241] = -18'sd     14;
assign PRECOMP_N1[242] = -18'sd     12;
assign PRECOMP_N1[243] = -18'sd      1;
assign PRECOMP_N1[244] =  18'sd     10;
assign PRECOMP_N1[245] =  18'sd     13;
assign PRECOMP_N1[246] =  18'sd      7;
assign PRECOMP_N1[247] = -18'sd      3;
assign PRECOMP_N1[248] = -18'sd     11;
assign PRECOMP_N1[249] = -18'sd     11;
assign PRECOMP_N1[250] = -18'sd      3;
assign PRECOMP_N1[251] =  18'sd      6;
assign PRECOMP_N1[252] =  18'sd     11;
assign PRECOMP_N1[253] =  18'sd      7;
assign PRECOMP_N1[254] = -18'sd      1;
assign PRECOMP_N1[255] = -18'sd      8;
assign PRECOMP_N1[256] = -18'sd      9;
assign PRECOMP_N1[257] = -18'sd      3;
assign PRECOMP_N1[258] =  18'sd      4;
assign PRECOMP_N1[259] =  18'sd      8;
assign PRECOMP_N1[260] =  18'sd      6;
assign PRECOMP_N1[261] = -18'sd      1;
assign PRECOMP_N1[262] = -18'sd      7;
assign PRECOMP_N1[263] = -18'sd      7;
assign PRECOMP_N1[264] = -18'sd      3;
assign PRECOMP_N1[265] =  18'sd      4;
assign PRECOMP_N1[266] =  18'sd      7;
assign PRECOMP_N1[267] =  18'sd      6;
assign PRECOMP_N1[268] =  18'sd      0;
assign PRECOMP_N1[269] = -18'sd      6;
assign PRECOMP_N1[270] = -18'sd      7;
assign PRECOMP_N1[271] = -18'sd      4;
assign PRECOMP_N1[272] =  18'sd      3;
assign PRECOMP_N1[273] =  18'sd      7;
assign PRECOMP_N1[274] =  18'sd      6;
assign PRECOMP_N1[275] =  18'sd      1;
assign PRECOMP_N1[276] = -18'sd      4;
assign PRECOMP_N1[277] = -18'sd      7;
assign PRECOMP_N1[278] = -18'sd      4;
assign PRECOMP_N1[279] =  18'sd      1;
assign PRECOMP_N1[280] =  18'sd      5;
assign PRECOMP_N1[281] =  18'sd      6;
assign PRECOMP_N1[282] =  18'sd      2;
assign PRECOMP_N1[283] = -18'sd      3;
assign PRECOMP_N1[284] = -18'sd      6;
assign PRECOMP_N1[285] = -18'sd      4;
assign PRECOMP_N1[286] =  18'sd      0;
assign PRECOMP_N1[287] =  18'sd      4;
assign PRECOMP_N1[288] =  18'sd      5;
assign PRECOMP_N1[289] =  18'sd      2;
assign PRECOMP_N1[290] = -18'sd      2;
assign PRECOMP_N1[291] = -18'sd      5;
assign PRECOMP_N1[292] = -18'sd      4;
assign PRECOMP_N1[293] =  18'sd      0;
assign PRECOMP_N1[294] =  18'sd      3;
assign PRECOMP_N1[295] =  18'sd      4;
assign PRECOMP_N1[296] =  18'sd      2;
assign PRECOMP_N1[297] = -18'sd      1;
assign PRECOMP_N1[298] = -18'sd      4;
assign PRECOMP_N1[299] = -18'sd      4;
assign PRECOMP_N1[300] = -18'sd      1;
assign PRECOMP_N1[301] =  18'sd      3;
assign PRECOMP_N1[302] =  18'sd      4;
assign PRECOMP_N1[303] =  18'sd      2;
assign PRECOMP_N1[304] = -18'sd      1;



//TX Filter 18'sd N2 LUT Coefficients (headroom)
assign PRECOMP_N2[  0] = -18'sd      3;
assign PRECOMP_N2[  1] =  18'sd      7;
assign PRECOMP_N2[  2] =  18'sd     12;
assign PRECOMP_N2[  3] =  18'sd      8;
assign PRECOMP_N2[  4] = -18'sd      2;
assign PRECOMP_N2[  5] = -18'sd     11;
assign PRECOMP_N2[  6] = -18'sd     12;
assign PRECOMP_N2[  7] = -18'sd      4;
assign PRECOMP_N2[  8] =  18'sd      7;
assign PRECOMP_N2[  9] =  18'sd     13;
assign PRECOMP_N2[ 10] =  18'sd     10;
assign PRECOMP_N2[ 11] = -18'sd      1;
assign PRECOMP_N2[ 12] = -18'sd     11;
assign PRECOMP_N2[ 13] = -18'sd     14;
assign PRECOMP_N2[ 14] = -18'sd      6;
assign PRECOMP_N2[ 15] =  18'sd      7;
assign PRECOMP_N2[ 16] =  18'sd     15;
assign PRECOMP_N2[ 17] =  18'sd     12;
assign PRECOMP_N2[ 18] =  18'sd      0;
assign PRECOMP_N2[ 19] = -18'sd     13;
assign PRECOMP_N2[ 20] = -18'sd     17;
assign PRECOMP_N2[ 21] = -18'sd      9;
assign PRECOMP_N2[ 22] =  18'sd      6;
assign PRECOMP_N2[ 23] =  18'sd     18;
assign PRECOMP_N2[ 24] =  18'sd     16;
assign PRECOMP_N2[ 25] =  18'sd      3;
assign PRECOMP_N2[ 26] = -18'sd     13;
assign PRECOMP_N2[ 27] = -18'sd     20;
assign PRECOMP_N2[ 28] = -18'sd     13;
assign PRECOMP_N2[ 29] =  18'sd      3;
assign PRECOMP_N2[ 30] =  18'sd     18;
assign PRECOMP_N2[ 31] =  18'sd     20;
assign PRECOMP_N2[ 32] =  18'sd      8;
assign PRECOMP_N2[ 33] = -18'sd     11;
assign PRECOMP_N2[ 34] = -18'sd     22;
assign PRECOMP_N2[ 35] = -18'sd     17;
assign PRECOMP_N2[ 36] =  18'sd      0;
assign PRECOMP_N2[ 37] =  18'sd     17;
assign PRECOMP_N2[ 38] =  18'sd     22;
assign PRECOMP_N2[ 39] =  18'sd     11;
assign PRECOMP_N2[ 40] = -18'sd      9;
assign PRECOMP_N2[ 41] = -18'sd     22;
assign PRECOMP_N2[ 42] = -18'sd     20;
assign PRECOMP_N2[ 43] = -18'sd      2;
assign PRECOMP_N2[ 44] =  18'sd     18;
assign PRECOMP_N2[ 45] =  18'sd     25;
assign PRECOMP_N2[ 46] =  18'sd     13;
assign PRECOMP_N2[ 47] = -18'sd      9;
assign PRECOMP_N2[ 48] = -18'sd     26;
assign PRECOMP_N2[ 49] = -18'sd     24;
assign PRECOMP_N2[ 50] = -18'sd      3;
assign PRECOMP_N2[ 51] =  18'sd     21;
assign PRECOMP_N2[ 52] =  18'sd     32;
assign PRECOMP_N2[ 53] =  18'sd     19;
assign PRECOMP_N2[ 54] = -18'sd      9;
assign PRECOMP_N2[ 55] = -18'sd     32;
assign PRECOMP_N2[ 56] = -18'sd     33;
assign PRECOMP_N2[ 57] = -18'sd     10;
assign PRECOMP_N2[ 58] =  18'sd     22;
assign PRECOMP_N2[ 59] =  18'sd     40;
assign PRECOMP_N2[ 60] =  18'sd     30;
assign PRECOMP_N2[ 61] = -18'sd      2;
assign PRECOMP_N2[ 62] = -18'sd     34;
assign PRECOMP_N2[ 63] = -18'sd     43;
assign PRECOMP_N2[ 64] = -18'sd     21;
assign PRECOMP_N2[ 65] =  18'sd     17;
assign PRECOMP_N2[ 66] =  18'sd     44;
assign PRECOMP_N2[ 67] =  18'sd     40;
assign PRECOMP_N2[ 68] =  18'sd      8;
assign PRECOMP_N2[ 69] = -18'sd     31;
assign PRECOMP_N2[ 70] = -18'sd     48;
assign PRECOMP_N2[ 71] = -18'sd     30;
assign PRECOMP_N2[ 72] =  18'sd     11;
assign PRECOMP_N2[ 73] =  18'sd     44;
assign PRECOMP_N2[ 74] =  18'sd     45;
assign PRECOMP_N2[ 75] =  18'sd     12;
assign PRECOMP_N2[ 76] = -18'sd     32;
assign PRECOMP_N2[ 77] = -18'sd     53;
assign PRECOMP_N2[ 78] = -18'sd     34;
assign PRECOMP_N2[ 79] =  18'sd     13;
assign PRECOMP_N2[ 80] =  18'sd     53;
assign PRECOMP_N2[ 81] =  18'sd     55;
assign PRECOMP_N2[ 82] =  18'sd     13;
assign PRECOMP_N2[ 83] = -18'sd     42;
assign PRECOMP_N2[ 84] = -18'sd     71;
assign PRECOMP_N2[ 85] = -18'sd     48;
assign PRECOMP_N2[ 86] =  18'sd     15;
assign PRECOMP_N2[ 87] =  18'sd     73;
assign PRECOMP_N2[ 88] =  18'sd     83;
assign PRECOMP_N2[ 89] =  18'sd     32;
assign PRECOMP_N2[ 90] = -18'sd     48;
assign PRECOMP_N2[ 91] = -18'sd    101;
assign PRECOMP_N2[ 92] = -18'sd     85;
assign PRECOMP_N2[ 93] = -18'sd      5;
assign PRECOMP_N2[ 94] =  18'sd     84;
assign PRECOMP_N2[ 95] =  18'sd    120;
assign PRECOMP_N2[ 96] =  18'sd     73;
assign PRECOMP_N2[ 97] = -18'sd     30;
assign PRECOMP_N2[ 98] = -18'sd    117;
assign PRECOMP_N2[ 99] = -18'sd    125;
assign PRECOMP_N2[100] = -18'sd     44;
assign PRECOMP_N2[101] =  18'sd     71;
assign PRECOMP_N2[102] =  18'sd    139;
assign PRECOMP_N2[103] =  18'sd    108;
assign PRECOMP_N2[104] = -18'sd      3;
assign PRECOMP_N2[105] = -18'sd    114;
assign PRECOMP_N2[106] = -18'sd    143;
assign PRECOMP_N2[107] = -18'sd     64;
assign PRECOMP_N2[108] =  18'sd     69;
assign PRECOMP_N2[109] =  18'sd    153;
assign PRECOMP_N2[110] =  18'sd    119;
assign PRECOMP_N2[111] = -18'sd     16;
assign PRECOMP_N2[112] = -18'sd    153;
assign PRECOMP_N2[113] = -18'sd    179;
assign PRECOMP_N2[114] = -18'sd     57;
assign PRECOMP_N2[115] =  18'sd    137;
assign PRECOMP_N2[116] =  18'sd    255;
assign PRECOMP_N2[117] =  18'sd    183;
assign PRECOMP_N2[118] = -18'sd     57;
assign PRECOMP_N2[119] = -18'sd    308;
assign PRECOMP_N2[120] = -18'sd    369;
assign PRECOMP_N2[121] = -18'sd    151;
assign PRECOMP_N2[122] =  18'sd    237;
assign PRECOMP_N2[123] =  18'sd    534;
assign PRECOMP_N2[124] =  18'sd    492;
assign PRECOMP_N2[125] =  18'sd     68;
assign PRECOMP_N2[126] = -18'sd    503;
assign PRECOMP_N2[127] = -18'sd    828;
assign PRECOMP_N2[128] = -18'sd    617;
assign PRECOMP_N2[129] =  18'sd     90;
assign PRECOMP_N2[130] =  18'sd    882;
assign PRECOMP_N2[131] =  18'sd   1208;
assign PRECOMP_N2[132] =  18'sd    738;
assign PRECOMP_N2[133] = -18'sd    357;
assign PRECOMP_N2[134] = -18'sd   1427;
assign PRECOMP_N2[135] = -18'sd   1713;
assign PRECOMP_N2[136] = -18'sd    848;
assign PRECOMP_N2[137] =  18'sd    801;
assign PRECOMP_N2[138] =  18'sd   2246;
assign PRECOMP_N2[139] =  18'sd   2432;
assign PRECOMP_N2[140] =  18'sd    942;
assign PRECOMP_N2[141] = -18'sd   1579;
assign PRECOMP_N2[142] = -18'sd   3622;
assign PRECOMP_N2[143] = -18'sd   3629;
assign PRECOMP_N2[144] = -18'sd   1013;
assign PRECOMP_N2[145] =  18'sd   3207;
assign PRECOMP_N2[146] =  18'sd   6607;
assign PRECOMP_N2[147] =  18'sd   6434;
assign PRECOMP_N2[148] =  18'sd   1057;
assign PRECOMP_N2[149] = -18'sd   8945;
assign PRECOMP_N2[150] = -18'sd  20712;
assign PRECOMP_N2[151] = -18'sd  30169;
assign PRECOMP_N2[152] = -18'sd  33785;
assign PRECOMP_N2[153] = -18'sd  30169;
assign PRECOMP_N2[154] = -18'sd  20712;
assign PRECOMP_N2[155] = -18'sd   8945;
assign PRECOMP_N2[156] =  18'sd   1057;
assign PRECOMP_N2[157] =  18'sd   6434;
assign PRECOMP_N2[158] =  18'sd   6607;
assign PRECOMP_N2[159] =  18'sd   3207;
assign PRECOMP_N2[160] = -18'sd   1013;
assign PRECOMP_N2[161] = -18'sd   3629;
assign PRECOMP_N2[162] = -18'sd   3622;
assign PRECOMP_N2[163] = -18'sd   1579;
assign PRECOMP_N2[164] =  18'sd    942;
assign PRECOMP_N2[165] =  18'sd   2432;
assign PRECOMP_N2[166] =  18'sd   2246;
assign PRECOMP_N2[167] =  18'sd    801;
assign PRECOMP_N2[168] = -18'sd    848;
assign PRECOMP_N2[169] = -18'sd   1713;
assign PRECOMP_N2[170] = -18'sd   1427;
assign PRECOMP_N2[171] = -18'sd    357;
assign PRECOMP_N2[172] =  18'sd    738;
assign PRECOMP_N2[173] =  18'sd   1208;
assign PRECOMP_N2[174] =  18'sd    882;
assign PRECOMP_N2[175] =  18'sd     90;
assign PRECOMP_N2[176] = -18'sd    617;
assign PRECOMP_N2[177] = -18'sd    828;
assign PRECOMP_N2[178] = -18'sd    503;
assign PRECOMP_N2[179] =  18'sd     68;
assign PRECOMP_N2[180] =  18'sd    492;
assign PRECOMP_N2[181] =  18'sd    534;
assign PRECOMP_N2[182] =  18'sd    237;
assign PRECOMP_N2[183] = -18'sd    151;
assign PRECOMP_N2[184] = -18'sd    369;
assign PRECOMP_N2[185] = -18'sd    308;
assign PRECOMP_N2[186] = -18'sd     57;
assign PRECOMP_N2[187] =  18'sd    183;
assign PRECOMP_N2[188] =  18'sd    255;
assign PRECOMP_N2[189] =  18'sd    137;
assign PRECOMP_N2[190] = -18'sd     57;
assign PRECOMP_N2[191] = -18'sd    179;
assign PRECOMP_N2[192] = -18'sd    153;
assign PRECOMP_N2[193] = -18'sd     16;
assign PRECOMP_N2[194] =  18'sd    119;
assign PRECOMP_N2[195] =  18'sd    153;
assign PRECOMP_N2[196] =  18'sd     69;
assign PRECOMP_N2[197] = -18'sd     64;
assign PRECOMP_N2[198] = -18'sd    143;
assign PRECOMP_N2[199] = -18'sd    114;
assign PRECOMP_N2[200] = -18'sd      3;
assign PRECOMP_N2[201] =  18'sd    108;
assign PRECOMP_N2[202] =  18'sd    139;
assign PRECOMP_N2[203] =  18'sd     71;
assign PRECOMP_N2[204] = -18'sd     44;
assign PRECOMP_N2[205] = -18'sd    125;
assign PRECOMP_N2[206] = -18'sd    117;
assign PRECOMP_N2[207] = -18'sd     30;
assign PRECOMP_N2[208] =  18'sd     73;
assign PRECOMP_N2[209] =  18'sd    120;
assign PRECOMP_N2[210] =  18'sd     84;
assign PRECOMP_N2[211] = -18'sd      5;
assign PRECOMP_N2[212] = -18'sd     85;
assign PRECOMP_N2[213] = -18'sd    101;
assign PRECOMP_N2[214] = -18'sd     48;
assign PRECOMP_N2[215] =  18'sd     32;
assign PRECOMP_N2[216] =  18'sd     83;
assign PRECOMP_N2[217] =  18'sd     73;
assign PRECOMP_N2[218] =  18'sd     15;
assign PRECOMP_N2[219] = -18'sd     48;
assign PRECOMP_N2[220] = -18'sd     71;
assign PRECOMP_N2[221] = -18'sd     42;
assign PRECOMP_N2[222] =  18'sd     13;
assign PRECOMP_N2[223] =  18'sd     55;
assign PRECOMP_N2[224] =  18'sd     53;
assign PRECOMP_N2[225] =  18'sd     13;
assign PRECOMP_N2[226] = -18'sd     34;
assign PRECOMP_N2[227] = -18'sd     53;
assign PRECOMP_N2[228] = -18'sd     32;
assign PRECOMP_N2[229] =  18'sd     12;
assign PRECOMP_N2[230] =  18'sd     45;
assign PRECOMP_N2[231] =  18'sd     44;
assign PRECOMP_N2[232] =  18'sd     11;
assign PRECOMP_N2[233] = -18'sd     30;
assign PRECOMP_N2[234] = -18'sd     48;
assign PRECOMP_N2[235] = -18'sd     31;
assign PRECOMP_N2[236] =  18'sd      8;
assign PRECOMP_N2[237] =  18'sd     40;
assign PRECOMP_N2[238] =  18'sd     44;
assign PRECOMP_N2[239] =  18'sd     17;
assign PRECOMP_N2[240] = -18'sd     21;
assign PRECOMP_N2[241] = -18'sd     43;
assign PRECOMP_N2[242] = -18'sd     34;
assign PRECOMP_N2[243] = -18'sd      2;
assign PRECOMP_N2[244] =  18'sd     30;
assign PRECOMP_N2[245] =  18'sd     40;
assign PRECOMP_N2[246] =  18'sd     22;
assign PRECOMP_N2[247] = -18'sd     10;
assign PRECOMP_N2[248] = -18'sd     33;
assign PRECOMP_N2[249] = -18'sd     32;
assign PRECOMP_N2[250] = -18'sd      9;
assign PRECOMP_N2[251] =  18'sd     19;
assign PRECOMP_N2[252] =  18'sd     32;
assign PRECOMP_N2[253] =  18'sd     21;
assign PRECOMP_N2[254] = -18'sd      3;
assign PRECOMP_N2[255] = -18'sd     24;
assign PRECOMP_N2[256] = -18'sd     26;
assign PRECOMP_N2[257] = -18'sd      9;
assign PRECOMP_N2[258] =  18'sd     13;
assign PRECOMP_N2[259] =  18'sd     25;
assign PRECOMP_N2[260] =  18'sd     18;
assign PRECOMP_N2[261] = -18'sd      2;
assign PRECOMP_N2[262] = -18'sd     20;
assign PRECOMP_N2[263] = -18'sd     22;
assign PRECOMP_N2[264] = -18'sd      9;
assign PRECOMP_N2[265] =  18'sd     11;
assign PRECOMP_N2[266] =  18'sd     22;
assign PRECOMP_N2[267] =  18'sd     17;
assign PRECOMP_N2[268] =  18'sd      0;
assign PRECOMP_N2[269] = -18'sd     17;
assign PRECOMP_N2[270] = -18'sd     22;
assign PRECOMP_N2[271] = -18'sd     11;
assign PRECOMP_N2[272] =  18'sd      8;
assign PRECOMP_N2[273] =  18'sd     20;
assign PRECOMP_N2[274] =  18'sd     18;
assign PRECOMP_N2[275] =  18'sd      3;
assign PRECOMP_N2[276] = -18'sd     13;
assign PRECOMP_N2[277] = -18'sd     20;
assign PRECOMP_N2[278] = -18'sd     13;
assign PRECOMP_N2[279] =  18'sd      3;
assign PRECOMP_N2[280] =  18'sd     16;
assign PRECOMP_N2[281] =  18'sd     18;
assign PRECOMP_N2[282] =  18'sd      6;
assign PRECOMP_N2[283] = -18'sd      9;
assign PRECOMP_N2[284] = -18'sd     17;
assign PRECOMP_N2[285] = -18'sd     13;
assign PRECOMP_N2[286] =  18'sd      0;
assign PRECOMP_N2[287] =  18'sd     12;
assign PRECOMP_N2[288] =  18'sd     15;
assign PRECOMP_N2[289] =  18'sd      7;
assign PRECOMP_N2[290] = -18'sd      6;
assign PRECOMP_N2[291] = -18'sd     14;
assign PRECOMP_N2[292] = -18'sd     11;
assign PRECOMP_N2[293] = -18'sd      1;
assign PRECOMP_N2[294] =  18'sd     10;
assign PRECOMP_N2[295] =  18'sd     13;
assign PRECOMP_N2[296] =  18'sd      7;
assign PRECOMP_N2[297] = -18'sd      4;
assign PRECOMP_N2[298] = -18'sd     12;
assign PRECOMP_N2[299] = -18'sd     11;
assign PRECOMP_N2[300] = -18'sd      2;
assign PRECOMP_N2[301] =  18'sd      8;
assign PRECOMP_N2[302] =  18'sd     12;
assign PRECOMP_N2[303] =  18'sd      7;
assign PRECOMP_N2[304] = -18'sd      3;


