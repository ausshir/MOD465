
//TX Filter 18'sd P2 LUT Coefficients (headroom)
assign PRECOMP_P2[  0] = -18'sd     24;
assign PRECOMP_P2[  1] = -18'sd      8;
assign PRECOMP_P2[  2] =  18'sd     15;
assign PRECOMP_P2[  3] =  18'sd     28;
assign PRECOMP_P2[  4] =  18'sd     21;
assign PRECOMP_P2[  5] = -18'sd      3;
assign PRECOMP_P2[  6] = -18'sd     26;
assign PRECOMP_P2[  7] = -18'sd     32;
assign PRECOMP_P2[  8] = -18'sd     13;
assign PRECOMP_P2[  9] =  18'sd     17;
assign PRECOMP_P2[ 10] =  18'sd     37;
assign PRECOMP_P2[ 11] =  18'sd     31;
assign PRECOMP_P2[ 12] =  18'sd      2;
assign PRECOMP_P2[ 13] = -18'sd     33;
assign PRECOMP_P2[ 14] = -18'sd     47;
assign PRECOMP_P2[ 15] = -18'sd     27;
assign PRECOMP_P2[ 16] =  18'sd     14;
assign PRECOMP_P2[ 17] =  18'sd     50;
assign PRECOMP_P2[ 18] =  18'sd     53;
assign PRECOMP_P2[ 19] =  18'sd     18;
assign PRECOMP_P2[ 20] = -18'sd     33;
assign PRECOMP_P2[ 21] = -18'sd     66;
assign PRECOMP_P2[ 22] = -18'sd     55;
assign PRECOMP_P2[ 23] = -18'sd      4;
assign PRECOMP_P2[ 24] =  18'sd     54;
assign PRECOMP_P2[ 25] =  18'sd     79;
assign PRECOMP_P2[ 26] =  18'sd     51;
assign PRECOMP_P2[ 27] = -18'sd     15;
assign PRECOMP_P2[ 28] = -18'sd     74;
assign PRECOMP_P2[ 29] = -18'sd     86;
assign PRECOMP_P2[ 30] = -18'sd     38;
assign PRECOMP_P2[ 31] =  18'sd     38;
assign PRECOMP_P2[ 32] =  18'sd     92;
assign PRECOMP_P2[ 33] =  18'sd     84;
assign PRECOMP_P2[ 34] =  18'sd     16;
assign PRECOMP_P2[ 35] = -18'sd     65;
assign PRECOMP_P2[ 36] = -18'sd    103;
assign PRECOMP_P2[ 37] = -18'sd     68;
assign PRECOMP_P2[ 38] =  18'sd     16;
assign PRECOMP_P2[ 39] =  18'sd     92;
assign PRECOMP_P2[ 40] =  18'sd    102;
assign PRECOMP_P2[ 41] =  18'sd     37;
assign PRECOMP_P2[ 42] = -18'sd     60;
assign PRECOMP_P2[ 43] = -18'sd    117;
assign PRECOMP_P2[ 44] = -18'sd     86;
assign PRECOMP_P2[ 45] =  18'sd     15;
assign PRECOMP_P2[ 46] =  18'sd    115;
assign PRECOMP_P2[ 47] =  18'sd    135;
assign PRECOMP_P2[ 48] =  18'sd     48;
assign PRECOMP_P2[ 49] = -18'sd     91;
assign PRECOMP_P2[ 50] = -18'sd    181;
assign PRECOMP_P2[ 51] = -18'sd    142;
assign PRECOMP_P2[ 52] =  18'sd     18;
assign PRECOMP_P2[ 53] =  18'sd    195;
assign PRECOMP_P2[ 54] =  18'sd    256;
assign PRECOMP_P2[ 55] =  18'sd    131;
assign PRECOMP_P2[ 56] = -18'sd    120;
assign PRECOMP_P2[ 57] = -18'sd    331;
assign PRECOMP_P2[ 58] = -18'sd    338;
assign PRECOMP_P2[ 59] = -18'sd     95;
assign PRECOMP_P2[ 60] =  18'sd    266;
assign PRECOMP_P2[ 61] =  18'sd    504;
assign PRECOMP_P2[ 62] =  18'sd    424;
assign PRECOMP_P2[ 63] =  18'sd     24;
assign PRECOMP_P2[ 64] = -18'sd    469;
assign PRECOMP_P2[ 65] = -18'sd    722;
assign PRECOMP_P2[ 66] = -18'sd    513;
assign PRECOMP_P2[ 67] =  18'sd     94;
assign PRECOMP_P2[ 68] =  18'sd    744;
assign PRECOMP_P2[ 69] =  18'sd    993;
assign PRECOMP_P2[ 70] =  18'sd    599;
assign PRECOMP_P2[ 71] = -18'sd    279;
assign PRECOMP_P2[ 72] = -18'sd   1120;
assign PRECOMP_P2[ 73] = -18'sd   1340;
assign PRECOMP_P2[ 74] = -18'sd    680;
assign PRECOMP_P2[ 75] =  18'sd    564;
assign PRECOMP_P2[ 76] =  18'sd   1647;
assign PRECOMP_P2[ 77] =  18'sd   1801;
assign PRECOMP_P2[ 78] =  18'sd    752;
assign PRECOMP_P2[ 79] = -18'sd   1014;
assign PRECOMP_P2[ 80] = -18'sd   2433;
assign PRECOMP_P2[ 81] = -18'sd   2471;
assign PRECOMP_P2[ 82] = -18'sd    811;
assign PRECOMP_P2[ 83] =  18'sd   1786;
assign PRECOMP_P2[ 84] =  18'sd   3765;
assign PRECOMP_P2[ 85] =  18'sd   3614;
assign PRECOMP_P2[ 86] =  18'sd    856;
assign PRECOMP_P2[ 87] = -18'sd   3393;
assign PRECOMP_P2[ 88] = -18'sd   6694;
assign PRECOMP_P2[ 89] = -18'sd   6364;
assign PRECOMP_P2[ 90] = -18'sd    884;
assign PRECOMP_P2[ 91] =  18'sd   9097;
assign PRECOMP_P2[ 92] =  18'sd  20733;
assign PRECOMP_P2[ 93] =  18'sd  30039;
assign PRECOMP_P2[ 94] =  18'sd  33589;
assign PRECOMP_P2[ 95] =  18'sd  30039;
assign PRECOMP_P2[ 96] =  18'sd  20733;
assign PRECOMP_P2[ 97] =  18'sd   9097;
assign PRECOMP_P2[ 98] = -18'sd    884;
assign PRECOMP_P2[ 99] = -18'sd   6364;
assign PRECOMP_P2[100] = -18'sd   6694;
assign PRECOMP_P2[101] = -18'sd   3393;
assign PRECOMP_P2[102] =  18'sd    856;
assign PRECOMP_P2[103] =  18'sd   3614;
assign PRECOMP_P2[104] =  18'sd   3765;
assign PRECOMP_P2[105] =  18'sd   1786;
assign PRECOMP_P2[106] = -18'sd    811;
assign PRECOMP_P2[107] = -18'sd   2471;
assign PRECOMP_P2[108] = -18'sd   2433;
assign PRECOMP_P2[109] = -18'sd   1014;
assign PRECOMP_P2[110] =  18'sd    752;
assign PRECOMP_P2[111] =  18'sd   1801;
assign PRECOMP_P2[112] =  18'sd   1647;
assign PRECOMP_P2[113] =  18'sd    564;
assign PRECOMP_P2[114] = -18'sd    680;
assign PRECOMP_P2[115] = -18'sd   1340;
assign PRECOMP_P2[116] = -18'sd   1120;
assign PRECOMP_P2[117] = -18'sd    279;
assign PRECOMP_P2[118] =  18'sd    599;
assign PRECOMP_P2[119] =  18'sd    993;
assign PRECOMP_P2[120] =  18'sd    744;
assign PRECOMP_P2[121] =  18'sd     94;
assign PRECOMP_P2[122] = -18'sd    513;
assign PRECOMP_P2[123] = -18'sd    722;
assign PRECOMP_P2[124] = -18'sd    469;
assign PRECOMP_P2[125] =  18'sd     24;
assign PRECOMP_P2[126] =  18'sd    424;
assign PRECOMP_P2[127] =  18'sd    504;
assign PRECOMP_P2[128] =  18'sd    266;
assign PRECOMP_P2[129] = -18'sd     95;
assign PRECOMP_P2[130] = -18'sd    338;
assign PRECOMP_P2[131] = -18'sd    331;
assign PRECOMP_P2[132] = -18'sd    120;
assign PRECOMP_P2[133] =  18'sd    131;
assign PRECOMP_P2[134] =  18'sd    256;
assign PRECOMP_P2[135] =  18'sd    195;
assign PRECOMP_P2[136] =  18'sd     18;
assign PRECOMP_P2[137] = -18'sd    142;
assign PRECOMP_P2[138] = -18'sd    181;
assign PRECOMP_P2[139] = -18'sd     91;
assign PRECOMP_P2[140] =  18'sd     48;
assign PRECOMP_P2[141] =  18'sd    135;
assign PRECOMP_P2[142] =  18'sd    115;
assign PRECOMP_P2[143] =  18'sd     15;
assign PRECOMP_P2[144] = -18'sd     86;
assign PRECOMP_P2[145] = -18'sd    117;
assign PRECOMP_P2[146] = -18'sd     60;
assign PRECOMP_P2[147] =  18'sd     37;
assign PRECOMP_P2[148] =  18'sd    102;
assign PRECOMP_P2[149] =  18'sd     92;
assign PRECOMP_P2[150] =  18'sd     16;
assign PRECOMP_P2[151] = -18'sd     68;
assign PRECOMP_P2[152] = -18'sd    103;
assign PRECOMP_P2[153] = -18'sd     65;
assign PRECOMP_P2[154] =  18'sd     16;
assign PRECOMP_P2[155] =  18'sd     84;
assign PRECOMP_P2[156] =  18'sd     92;
assign PRECOMP_P2[157] =  18'sd     38;
assign PRECOMP_P2[158] = -18'sd     38;
assign PRECOMP_P2[159] = -18'sd     86;
assign PRECOMP_P2[160] = -18'sd     74;
assign PRECOMP_P2[161] = -18'sd     15;
assign PRECOMP_P2[162] =  18'sd     51;
assign PRECOMP_P2[163] =  18'sd     79;
assign PRECOMP_P2[164] =  18'sd     54;
assign PRECOMP_P2[165] = -18'sd      4;
assign PRECOMP_P2[166] = -18'sd     55;
assign PRECOMP_P2[167] = -18'sd     66;
assign PRECOMP_P2[168] = -18'sd     33;
assign PRECOMP_P2[169] =  18'sd     18;
assign PRECOMP_P2[170] =  18'sd     53;
assign PRECOMP_P2[171] =  18'sd     50;
assign PRECOMP_P2[172] =  18'sd     14;
assign PRECOMP_P2[173] = -18'sd     27;
assign PRECOMP_P2[174] = -18'sd     47;
assign PRECOMP_P2[175] = -18'sd     33;
assign PRECOMP_P2[176] =  18'sd      2;
assign PRECOMP_P2[177] =  18'sd     31;
assign PRECOMP_P2[178] =  18'sd     37;
assign PRECOMP_P2[179] =  18'sd     17;
assign PRECOMP_P2[180] = -18'sd     13;
assign PRECOMP_P2[181] = -18'sd     32;
assign PRECOMP_P2[182] = -18'sd     26;
assign PRECOMP_P2[183] = -18'sd      3;
assign PRECOMP_P2[184] =  18'sd     21;
assign PRECOMP_P2[185] =  18'sd     28;
assign PRECOMP_P2[186] =  18'sd     15;
assign PRECOMP_P2[187] = -18'sd      8;
assign PRECOMP_P2[188] = -18'sd     24;



//TX Filter 18'sd P1 LUT Coefficients (headroom)
assign PRECOMP_P1[  0] = -18'sd      8;
assign PRECOMP_P1[  1] = -18'sd      3;
assign PRECOMP_P1[  2] =  18'sd      5;
assign PRECOMP_P1[  3] =  18'sd      9;
assign PRECOMP_P1[  4] =  18'sd      7;
assign PRECOMP_P1[  5] = -18'sd      1;
assign PRECOMP_P1[  6] = -18'sd      9;
assign PRECOMP_P1[  7] = -18'sd     11;
assign PRECOMP_P1[  8] = -18'sd      4;
assign PRECOMP_P1[  9] =  18'sd      6;
assign PRECOMP_P1[ 10] =  18'sd     12;
assign PRECOMP_P1[ 11] =  18'sd     11;
assign PRECOMP_P1[ 12] =  18'sd      1;
assign PRECOMP_P1[ 13] = -18'sd     11;
assign PRECOMP_P1[ 14] = -18'sd     16;
assign PRECOMP_P1[ 15] = -18'sd      9;
assign PRECOMP_P1[ 16] =  18'sd      5;
assign PRECOMP_P1[ 17] =  18'sd     17;
assign PRECOMP_P1[ 18] =  18'sd     18;
assign PRECOMP_P1[ 19] =  18'sd      6;
assign PRECOMP_P1[ 20] = -18'sd     11;
assign PRECOMP_P1[ 21] = -18'sd     22;
assign PRECOMP_P1[ 22] = -18'sd     18;
assign PRECOMP_P1[ 23] = -18'sd      1;
assign PRECOMP_P1[ 24] =  18'sd     18;
assign PRECOMP_P1[ 25] =  18'sd     26;
assign PRECOMP_P1[ 26] =  18'sd     17;
assign PRECOMP_P1[ 27] = -18'sd      5;
assign PRECOMP_P1[ 28] = -18'sd     25;
assign PRECOMP_P1[ 29] = -18'sd     29;
assign PRECOMP_P1[ 30] = -18'sd     13;
assign PRECOMP_P1[ 31] =  18'sd     13;
assign PRECOMP_P1[ 32] =  18'sd     31;
assign PRECOMP_P1[ 33] =  18'sd     28;
assign PRECOMP_P1[ 34] =  18'sd      5;
assign PRECOMP_P1[ 35] = -18'sd     22;
assign PRECOMP_P1[ 36] = -18'sd     34;
assign PRECOMP_P1[ 37] = -18'sd     23;
assign PRECOMP_P1[ 38] =  18'sd      5;
assign PRECOMP_P1[ 39] =  18'sd     31;
assign PRECOMP_P1[ 40] =  18'sd     34;
assign PRECOMP_P1[ 41] =  18'sd     12;
assign PRECOMP_P1[ 42] = -18'sd     20;
assign PRECOMP_P1[ 43] = -18'sd     39;
assign PRECOMP_P1[ 44] = -18'sd     29;
assign PRECOMP_P1[ 45] =  18'sd      5;
assign PRECOMP_P1[ 46] =  18'sd     38;
assign PRECOMP_P1[ 47] =  18'sd     45;
assign PRECOMP_P1[ 48] =  18'sd     16;
assign PRECOMP_P1[ 49] = -18'sd     30;
assign PRECOMP_P1[ 50] = -18'sd     60;
assign PRECOMP_P1[ 51] = -18'sd     47;
assign PRECOMP_P1[ 52] =  18'sd      6;
assign PRECOMP_P1[ 53] =  18'sd     65;
assign PRECOMP_P1[ 54] =  18'sd     85;
assign PRECOMP_P1[ 55] =  18'sd     44;
assign PRECOMP_P1[ 56] = -18'sd     40;
assign PRECOMP_P1[ 57] = -18'sd    111;
assign PRECOMP_P1[ 58] = -18'sd    113;
assign PRECOMP_P1[ 59] = -18'sd     32;
assign PRECOMP_P1[ 60] =  18'sd     89;
assign PRECOMP_P1[ 61] =  18'sd    168;
assign PRECOMP_P1[ 62] =  18'sd    142;
assign PRECOMP_P1[ 63] =  18'sd      8;
assign PRECOMP_P1[ 64] = -18'sd    156;
assign PRECOMP_P1[ 65] = -18'sd    241;
assign PRECOMP_P1[ 66] = -18'sd    171;
assign PRECOMP_P1[ 67] =  18'sd     31;
assign PRECOMP_P1[ 68] =  18'sd    249;
assign PRECOMP_P1[ 69] =  18'sd    332;
assign PRECOMP_P1[ 70] =  18'sd    200;
assign PRECOMP_P1[ 71] = -18'sd     93;
assign PRECOMP_P1[ 72] = -18'sd    374;
assign PRECOMP_P1[ 73] = -18'sd    448;
assign PRECOMP_P1[ 74] = -18'sd    227;
assign PRECOMP_P1[ 75] =  18'sd    188;
assign PRECOMP_P1[ 76] =  18'sd    550;
assign PRECOMP_P1[ 77] =  18'sd    602;
assign PRECOMP_P1[ 78] =  18'sd    251;
assign PRECOMP_P1[ 79] = -18'sd    339;
assign PRECOMP_P1[ 80] = -18'sd    813;
assign PRECOMP_P1[ 81] = -18'sd    825;
assign PRECOMP_P1[ 82] = -18'sd    271;
assign PRECOMP_P1[ 83] =  18'sd    596;
assign PRECOMP_P1[ 84] =  18'sd   1257;
assign PRECOMP_P1[ 85] =  18'sd   1207;
assign PRECOMP_P1[ 86] =  18'sd    286;
assign PRECOMP_P1[ 87] = -18'sd   1133;
assign PRECOMP_P1[ 88] = -18'sd   2236;
assign PRECOMP_P1[ 89] = -18'sd   2126;
assign PRECOMP_P1[ 90] = -18'sd    295;
assign PRECOMP_P1[ 91] =  18'sd   3038;
assign PRECOMP_P1[ 92] =  18'sd   6925;
assign PRECOMP_P1[ 93] =  18'sd  10033;
assign PRECOMP_P1[ 94] =  18'sd  11219;
assign PRECOMP_P1[ 95] =  18'sd  10033;
assign PRECOMP_P1[ 96] =  18'sd   6925;
assign PRECOMP_P1[ 97] =  18'sd   3038;
assign PRECOMP_P1[ 98] = -18'sd    295;
assign PRECOMP_P1[ 99] = -18'sd   2126;
assign PRECOMP_P1[100] = -18'sd   2236;
assign PRECOMP_P1[101] = -18'sd   1133;
assign PRECOMP_P1[102] =  18'sd    286;
assign PRECOMP_P1[103] =  18'sd   1207;
assign PRECOMP_P1[104] =  18'sd   1257;
assign PRECOMP_P1[105] =  18'sd    596;
assign PRECOMP_P1[106] = -18'sd    271;
assign PRECOMP_P1[107] = -18'sd    825;
assign PRECOMP_P1[108] = -18'sd    813;
assign PRECOMP_P1[109] = -18'sd    339;
assign PRECOMP_P1[110] =  18'sd    251;
assign PRECOMP_P1[111] =  18'sd    602;
assign PRECOMP_P1[112] =  18'sd    550;
assign PRECOMP_P1[113] =  18'sd    188;
assign PRECOMP_P1[114] = -18'sd    227;
assign PRECOMP_P1[115] = -18'sd    448;
assign PRECOMP_P1[116] = -18'sd    374;
assign PRECOMP_P1[117] = -18'sd     93;
assign PRECOMP_P1[118] =  18'sd    200;
assign PRECOMP_P1[119] =  18'sd    332;
assign PRECOMP_P1[120] =  18'sd    249;
assign PRECOMP_P1[121] =  18'sd     31;
assign PRECOMP_P1[122] = -18'sd    171;
assign PRECOMP_P1[123] = -18'sd    241;
assign PRECOMP_P1[124] = -18'sd    156;
assign PRECOMP_P1[125] =  18'sd      8;
assign PRECOMP_P1[126] =  18'sd    142;
assign PRECOMP_P1[127] =  18'sd    168;
assign PRECOMP_P1[128] =  18'sd     89;
assign PRECOMP_P1[129] = -18'sd     32;
assign PRECOMP_P1[130] = -18'sd    113;
assign PRECOMP_P1[131] = -18'sd    111;
assign PRECOMP_P1[132] = -18'sd     40;
assign PRECOMP_P1[133] =  18'sd     44;
assign PRECOMP_P1[134] =  18'sd     85;
assign PRECOMP_P1[135] =  18'sd     65;
assign PRECOMP_P1[136] =  18'sd      6;
assign PRECOMP_P1[137] = -18'sd     47;
assign PRECOMP_P1[138] = -18'sd     60;
assign PRECOMP_P1[139] = -18'sd     30;
assign PRECOMP_P1[140] =  18'sd     16;
assign PRECOMP_P1[141] =  18'sd     45;
assign PRECOMP_P1[142] =  18'sd     38;
assign PRECOMP_P1[143] =  18'sd      5;
assign PRECOMP_P1[144] = -18'sd     29;
assign PRECOMP_P1[145] = -18'sd     39;
assign PRECOMP_P1[146] = -18'sd     20;
assign PRECOMP_P1[147] =  18'sd     12;
assign PRECOMP_P1[148] =  18'sd     34;
assign PRECOMP_P1[149] =  18'sd     31;
assign PRECOMP_P1[150] =  18'sd      5;
assign PRECOMP_P1[151] = -18'sd     23;
assign PRECOMP_P1[152] = -18'sd     34;
assign PRECOMP_P1[153] = -18'sd     22;
assign PRECOMP_P1[154] =  18'sd      5;
assign PRECOMP_P1[155] =  18'sd     28;
assign PRECOMP_P1[156] =  18'sd     31;
assign PRECOMP_P1[157] =  18'sd     13;
assign PRECOMP_P1[158] = -18'sd     13;
assign PRECOMP_P1[159] = -18'sd     29;
assign PRECOMP_P1[160] = -18'sd     25;
assign PRECOMP_P1[161] = -18'sd      5;
assign PRECOMP_P1[162] =  18'sd     17;
assign PRECOMP_P1[163] =  18'sd     26;
assign PRECOMP_P1[164] =  18'sd     18;
assign PRECOMP_P1[165] = -18'sd      1;
assign PRECOMP_P1[166] = -18'sd     18;
assign PRECOMP_P1[167] = -18'sd     22;
assign PRECOMP_P1[168] = -18'sd     11;
assign PRECOMP_P1[169] =  18'sd      6;
assign PRECOMP_P1[170] =  18'sd     18;
assign PRECOMP_P1[171] =  18'sd     17;
assign PRECOMP_P1[172] =  18'sd      5;
assign PRECOMP_P1[173] = -18'sd      9;
assign PRECOMP_P1[174] = -18'sd     16;
assign PRECOMP_P1[175] = -18'sd     11;
assign PRECOMP_P1[176] =  18'sd      1;
assign PRECOMP_P1[177] =  18'sd     11;
assign PRECOMP_P1[178] =  18'sd     12;
assign PRECOMP_P1[179] =  18'sd      6;
assign PRECOMP_P1[180] = -18'sd      4;
assign PRECOMP_P1[181] = -18'sd     11;
assign PRECOMP_P1[182] = -18'sd      9;
assign PRECOMP_P1[183] = -18'sd      1;
assign PRECOMP_P1[184] =  18'sd      7;
assign PRECOMP_P1[185] =  18'sd      9;
assign PRECOMP_P1[186] =  18'sd      5;
assign PRECOMP_P1[187] = -18'sd      3;
assign PRECOMP_P1[188] = -18'sd      8;



//TX Filter 18'sd N1 LUT Coefficients (headroom)
assign PRECOMP_N1[  0] =  18'sd      8;
assign PRECOMP_N1[  1] =  18'sd      3;
assign PRECOMP_N1[  2] = -18'sd      5;
assign PRECOMP_N1[  3] = -18'sd      9;
assign PRECOMP_N1[  4] = -18'sd      7;
assign PRECOMP_N1[  5] =  18'sd      1;
assign PRECOMP_N1[  6] =  18'sd      9;
assign PRECOMP_N1[  7] =  18'sd     11;
assign PRECOMP_N1[  8] =  18'sd      4;
assign PRECOMP_N1[  9] = -18'sd      6;
assign PRECOMP_N1[ 10] = -18'sd     12;
assign PRECOMP_N1[ 11] = -18'sd     11;
assign PRECOMP_N1[ 12] = -18'sd      1;
assign PRECOMP_N1[ 13] =  18'sd     11;
assign PRECOMP_N1[ 14] =  18'sd     16;
assign PRECOMP_N1[ 15] =  18'sd      9;
assign PRECOMP_N1[ 16] = -18'sd      5;
assign PRECOMP_N1[ 17] = -18'sd     17;
assign PRECOMP_N1[ 18] = -18'sd     18;
assign PRECOMP_N1[ 19] = -18'sd      6;
assign PRECOMP_N1[ 20] =  18'sd     11;
assign PRECOMP_N1[ 21] =  18'sd     22;
assign PRECOMP_N1[ 22] =  18'sd     18;
assign PRECOMP_N1[ 23] =  18'sd      1;
assign PRECOMP_N1[ 24] = -18'sd     18;
assign PRECOMP_N1[ 25] = -18'sd     26;
assign PRECOMP_N1[ 26] = -18'sd     17;
assign PRECOMP_N1[ 27] =  18'sd      5;
assign PRECOMP_N1[ 28] =  18'sd     25;
assign PRECOMP_N1[ 29] =  18'sd     29;
assign PRECOMP_N1[ 30] =  18'sd     13;
assign PRECOMP_N1[ 31] = -18'sd     13;
assign PRECOMP_N1[ 32] = -18'sd     31;
assign PRECOMP_N1[ 33] = -18'sd     28;
assign PRECOMP_N1[ 34] = -18'sd      5;
assign PRECOMP_N1[ 35] =  18'sd     22;
assign PRECOMP_N1[ 36] =  18'sd     34;
assign PRECOMP_N1[ 37] =  18'sd     23;
assign PRECOMP_N1[ 38] = -18'sd      5;
assign PRECOMP_N1[ 39] = -18'sd     31;
assign PRECOMP_N1[ 40] = -18'sd     34;
assign PRECOMP_N1[ 41] = -18'sd     12;
assign PRECOMP_N1[ 42] =  18'sd     20;
assign PRECOMP_N1[ 43] =  18'sd     39;
assign PRECOMP_N1[ 44] =  18'sd     29;
assign PRECOMP_N1[ 45] = -18'sd      5;
assign PRECOMP_N1[ 46] = -18'sd     38;
assign PRECOMP_N1[ 47] = -18'sd     45;
assign PRECOMP_N1[ 48] = -18'sd     16;
assign PRECOMP_N1[ 49] =  18'sd     30;
assign PRECOMP_N1[ 50] =  18'sd     60;
assign PRECOMP_N1[ 51] =  18'sd     47;
assign PRECOMP_N1[ 52] = -18'sd      6;
assign PRECOMP_N1[ 53] = -18'sd     65;
assign PRECOMP_N1[ 54] = -18'sd     85;
assign PRECOMP_N1[ 55] = -18'sd     44;
assign PRECOMP_N1[ 56] =  18'sd     40;
assign PRECOMP_N1[ 57] =  18'sd    111;
assign PRECOMP_N1[ 58] =  18'sd    113;
assign PRECOMP_N1[ 59] =  18'sd     32;
assign PRECOMP_N1[ 60] = -18'sd     89;
assign PRECOMP_N1[ 61] = -18'sd    168;
assign PRECOMP_N1[ 62] = -18'sd    142;
assign PRECOMP_N1[ 63] = -18'sd      8;
assign PRECOMP_N1[ 64] =  18'sd    156;
assign PRECOMP_N1[ 65] =  18'sd    241;
assign PRECOMP_N1[ 66] =  18'sd    171;
assign PRECOMP_N1[ 67] = -18'sd     31;
assign PRECOMP_N1[ 68] = -18'sd    249;
assign PRECOMP_N1[ 69] = -18'sd    332;
assign PRECOMP_N1[ 70] = -18'sd    200;
assign PRECOMP_N1[ 71] =  18'sd     93;
assign PRECOMP_N1[ 72] =  18'sd    374;
assign PRECOMP_N1[ 73] =  18'sd    448;
assign PRECOMP_N1[ 74] =  18'sd    227;
assign PRECOMP_N1[ 75] = -18'sd    188;
assign PRECOMP_N1[ 76] = -18'sd    550;
assign PRECOMP_N1[ 77] = -18'sd    602;
assign PRECOMP_N1[ 78] = -18'sd    251;
assign PRECOMP_N1[ 79] =  18'sd    339;
assign PRECOMP_N1[ 80] =  18'sd    813;
assign PRECOMP_N1[ 81] =  18'sd    825;
assign PRECOMP_N1[ 82] =  18'sd    271;
assign PRECOMP_N1[ 83] = -18'sd    596;
assign PRECOMP_N1[ 84] = -18'sd   1257;
assign PRECOMP_N1[ 85] = -18'sd   1207;
assign PRECOMP_N1[ 86] = -18'sd    286;
assign PRECOMP_N1[ 87] =  18'sd   1133;
assign PRECOMP_N1[ 88] =  18'sd   2236;
assign PRECOMP_N1[ 89] =  18'sd   2126;
assign PRECOMP_N1[ 90] =  18'sd    295;
assign PRECOMP_N1[ 91] = -18'sd   3038;
assign PRECOMP_N1[ 92] = -18'sd   6925;
assign PRECOMP_N1[ 93] = -18'sd  10033;
assign PRECOMP_N1[ 94] = -18'sd  11219;
assign PRECOMP_N1[ 95] = -18'sd  10033;
assign PRECOMP_N1[ 96] = -18'sd   6925;
assign PRECOMP_N1[ 97] = -18'sd   3038;
assign PRECOMP_N1[ 98] =  18'sd    295;
assign PRECOMP_N1[ 99] =  18'sd   2126;
assign PRECOMP_N1[100] =  18'sd   2236;
assign PRECOMP_N1[101] =  18'sd   1133;
assign PRECOMP_N1[102] = -18'sd    286;
assign PRECOMP_N1[103] = -18'sd   1207;
assign PRECOMP_N1[104] = -18'sd   1257;
assign PRECOMP_N1[105] = -18'sd    596;
assign PRECOMP_N1[106] =  18'sd    271;
assign PRECOMP_N1[107] =  18'sd    825;
assign PRECOMP_N1[108] =  18'sd    813;
assign PRECOMP_N1[109] =  18'sd    339;
assign PRECOMP_N1[110] = -18'sd    251;
assign PRECOMP_N1[111] = -18'sd    602;
assign PRECOMP_N1[112] = -18'sd    550;
assign PRECOMP_N1[113] = -18'sd    188;
assign PRECOMP_N1[114] =  18'sd    227;
assign PRECOMP_N1[115] =  18'sd    448;
assign PRECOMP_N1[116] =  18'sd    374;
assign PRECOMP_N1[117] =  18'sd     93;
assign PRECOMP_N1[118] = -18'sd    200;
assign PRECOMP_N1[119] = -18'sd    332;
assign PRECOMP_N1[120] = -18'sd    249;
assign PRECOMP_N1[121] = -18'sd     31;
assign PRECOMP_N1[122] =  18'sd    171;
assign PRECOMP_N1[123] =  18'sd    241;
assign PRECOMP_N1[124] =  18'sd    156;
assign PRECOMP_N1[125] = -18'sd      8;
assign PRECOMP_N1[126] = -18'sd    142;
assign PRECOMP_N1[127] = -18'sd    168;
assign PRECOMP_N1[128] = -18'sd     89;
assign PRECOMP_N1[129] =  18'sd     32;
assign PRECOMP_N1[130] =  18'sd    113;
assign PRECOMP_N1[131] =  18'sd    111;
assign PRECOMP_N1[132] =  18'sd     40;
assign PRECOMP_N1[133] = -18'sd     44;
assign PRECOMP_N1[134] = -18'sd     85;
assign PRECOMP_N1[135] = -18'sd     65;
assign PRECOMP_N1[136] = -18'sd      6;
assign PRECOMP_N1[137] =  18'sd     47;
assign PRECOMP_N1[138] =  18'sd     60;
assign PRECOMP_N1[139] =  18'sd     30;
assign PRECOMP_N1[140] = -18'sd     16;
assign PRECOMP_N1[141] = -18'sd     45;
assign PRECOMP_N1[142] = -18'sd     38;
assign PRECOMP_N1[143] = -18'sd      5;
assign PRECOMP_N1[144] =  18'sd     29;
assign PRECOMP_N1[145] =  18'sd     39;
assign PRECOMP_N1[146] =  18'sd     20;
assign PRECOMP_N1[147] = -18'sd     12;
assign PRECOMP_N1[148] = -18'sd     34;
assign PRECOMP_N1[149] = -18'sd     31;
assign PRECOMP_N1[150] = -18'sd      5;
assign PRECOMP_N1[151] =  18'sd     23;
assign PRECOMP_N1[152] =  18'sd     34;
assign PRECOMP_N1[153] =  18'sd     22;
assign PRECOMP_N1[154] = -18'sd      5;
assign PRECOMP_N1[155] = -18'sd     28;
assign PRECOMP_N1[156] = -18'sd     31;
assign PRECOMP_N1[157] = -18'sd     13;
assign PRECOMP_N1[158] =  18'sd     13;
assign PRECOMP_N1[159] =  18'sd     29;
assign PRECOMP_N1[160] =  18'sd     25;
assign PRECOMP_N1[161] =  18'sd      5;
assign PRECOMP_N1[162] = -18'sd     17;
assign PRECOMP_N1[163] = -18'sd     26;
assign PRECOMP_N1[164] = -18'sd     18;
assign PRECOMP_N1[165] =  18'sd      1;
assign PRECOMP_N1[166] =  18'sd     18;
assign PRECOMP_N1[167] =  18'sd     22;
assign PRECOMP_N1[168] =  18'sd     11;
assign PRECOMP_N1[169] = -18'sd      6;
assign PRECOMP_N1[170] = -18'sd     18;
assign PRECOMP_N1[171] = -18'sd     17;
assign PRECOMP_N1[172] = -18'sd      5;
assign PRECOMP_N1[173] =  18'sd      9;
assign PRECOMP_N1[174] =  18'sd     16;
assign PRECOMP_N1[175] =  18'sd     11;
assign PRECOMP_N1[176] = -18'sd      1;
assign PRECOMP_N1[177] = -18'sd     11;
assign PRECOMP_N1[178] = -18'sd     12;
assign PRECOMP_N1[179] = -18'sd      6;
assign PRECOMP_N1[180] =  18'sd      4;
assign PRECOMP_N1[181] =  18'sd     11;
assign PRECOMP_N1[182] =  18'sd      9;
assign PRECOMP_N1[183] =  18'sd      1;
assign PRECOMP_N1[184] = -18'sd      7;
assign PRECOMP_N1[185] = -18'sd      9;
assign PRECOMP_N1[186] = -18'sd      5;
assign PRECOMP_N1[187] =  18'sd      3;
assign PRECOMP_N1[188] =  18'sd      8;



//TX Filter 18'sd N2 LUT Coefficients (headroom)
assign PRECOMP_N2[  0] =  18'sd     24;
assign PRECOMP_N2[  1] =  18'sd      8;
assign PRECOMP_N2[  2] = -18'sd     15;
assign PRECOMP_N2[  3] = -18'sd     28;
assign PRECOMP_N2[  4] = -18'sd     21;
assign PRECOMP_N2[  5] =  18'sd      3;
assign PRECOMP_N2[  6] =  18'sd     26;
assign PRECOMP_N2[  7] =  18'sd     32;
assign PRECOMP_N2[  8] =  18'sd     13;
assign PRECOMP_N2[  9] = -18'sd     17;
assign PRECOMP_N2[ 10] = -18'sd     37;
assign PRECOMP_N2[ 11] = -18'sd     31;
assign PRECOMP_N2[ 12] = -18'sd      2;
assign PRECOMP_N2[ 13] =  18'sd     33;
assign PRECOMP_N2[ 14] =  18'sd     47;
assign PRECOMP_N2[ 15] =  18'sd     27;
assign PRECOMP_N2[ 16] = -18'sd     14;
assign PRECOMP_N2[ 17] = -18'sd     50;
assign PRECOMP_N2[ 18] = -18'sd     53;
assign PRECOMP_N2[ 19] = -18'sd     18;
assign PRECOMP_N2[ 20] =  18'sd     33;
assign PRECOMP_N2[ 21] =  18'sd     66;
assign PRECOMP_N2[ 22] =  18'sd     55;
assign PRECOMP_N2[ 23] =  18'sd      4;
assign PRECOMP_N2[ 24] = -18'sd     54;
assign PRECOMP_N2[ 25] = -18'sd     79;
assign PRECOMP_N2[ 26] = -18'sd     51;
assign PRECOMP_N2[ 27] =  18'sd     15;
assign PRECOMP_N2[ 28] =  18'sd     74;
assign PRECOMP_N2[ 29] =  18'sd     86;
assign PRECOMP_N2[ 30] =  18'sd     38;
assign PRECOMP_N2[ 31] = -18'sd     38;
assign PRECOMP_N2[ 32] = -18'sd     92;
assign PRECOMP_N2[ 33] = -18'sd     84;
assign PRECOMP_N2[ 34] = -18'sd     16;
assign PRECOMP_N2[ 35] =  18'sd     65;
assign PRECOMP_N2[ 36] =  18'sd    103;
assign PRECOMP_N2[ 37] =  18'sd     68;
assign PRECOMP_N2[ 38] = -18'sd     16;
assign PRECOMP_N2[ 39] = -18'sd     92;
assign PRECOMP_N2[ 40] = -18'sd    102;
assign PRECOMP_N2[ 41] = -18'sd     37;
assign PRECOMP_N2[ 42] =  18'sd     60;
assign PRECOMP_N2[ 43] =  18'sd    117;
assign PRECOMP_N2[ 44] =  18'sd     86;
assign PRECOMP_N2[ 45] = -18'sd     15;
assign PRECOMP_N2[ 46] = -18'sd    115;
assign PRECOMP_N2[ 47] = -18'sd    135;
assign PRECOMP_N2[ 48] = -18'sd     48;
assign PRECOMP_N2[ 49] =  18'sd     91;
assign PRECOMP_N2[ 50] =  18'sd    181;
assign PRECOMP_N2[ 51] =  18'sd    142;
assign PRECOMP_N2[ 52] = -18'sd     18;
assign PRECOMP_N2[ 53] = -18'sd    195;
assign PRECOMP_N2[ 54] = -18'sd    256;
assign PRECOMP_N2[ 55] = -18'sd    131;
assign PRECOMP_N2[ 56] =  18'sd    120;
assign PRECOMP_N2[ 57] =  18'sd    331;
assign PRECOMP_N2[ 58] =  18'sd    338;
assign PRECOMP_N2[ 59] =  18'sd     95;
assign PRECOMP_N2[ 60] = -18'sd    266;
assign PRECOMP_N2[ 61] = -18'sd    504;
assign PRECOMP_N2[ 62] = -18'sd    424;
assign PRECOMP_N2[ 63] = -18'sd     24;
assign PRECOMP_N2[ 64] =  18'sd    469;
assign PRECOMP_N2[ 65] =  18'sd    722;
assign PRECOMP_N2[ 66] =  18'sd    513;
assign PRECOMP_N2[ 67] = -18'sd     94;
assign PRECOMP_N2[ 68] = -18'sd    744;
assign PRECOMP_N2[ 69] = -18'sd    993;
assign PRECOMP_N2[ 70] = -18'sd    599;
assign PRECOMP_N2[ 71] =  18'sd    279;
assign PRECOMP_N2[ 72] =  18'sd   1120;
assign PRECOMP_N2[ 73] =  18'sd   1340;
assign PRECOMP_N2[ 74] =  18'sd    680;
assign PRECOMP_N2[ 75] = -18'sd    564;
assign PRECOMP_N2[ 76] = -18'sd   1647;
assign PRECOMP_N2[ 77] = -18'sd   1801;
assign PRECOMP_N2[ 78] = -18'sd    752;
assign PRECOMP_N2[ 79] =  18'sd   1014;
assign PRECOMP_N2[ 80] =  18'sd   2433;
assign PRECOMP_N2[ 81] =  18'sd   2471;
assign PRECOMP_N2[ 82] =  18'sd    811;
assign PRECOMP_N2[ 83] = -18'sd   1786;
assign PRECOMP_N2[ 84] = -18'sd   3765;
assign PRECOMP_N2[ 85] = -18'sd   3614;
assign PRECOMP_N2[ 86] = -18'sd    856;
assign PRECOMP_N2[ 87] =  18'sd   3393;
assign PRECOMP_N2[ 88] =  18'sd   6694;
assign PRECOMP_N2[ 89] =  18'sd   6364;
assign PRECOMP_N2[ 90] =  18'sd    884;
assign PRECOMP_N2[ 91] = -18'sd   9097;
assign PRECOMP_N2[ 92] = -18'sd  20733;
assign PRECOMP_N2[ 93] = -18'sd  30039;
assign PRECOMP_N2[ 94] = -18'sd  33589;
assign PRECOMP_N2[ 95] = -18'sd  30039;
assign PRECOMP_N2[ 96] = -18'sd  20733;
assign PRECOMP_N2[ 97] = -18'sd   9097;
assign PRECOMP_N2[ 98] =  18'sd    884;
assign PRECOMP_N2[ 99] =  18'sd   6364;
assign PRECOMP_N2[100] =  18'sd   6694;
assign PRECOMP_N2[101] =  18'sd   3393;
assign PRECOMP_N2[102] = -18'sd    856;
assign PRECOMP_N2[103] = -18'sd   3614;
assign PRECOMP_N2[104] = -18'sd   3765;
assign PRECOMP_N2[105] = -18'sd   1786;
assign PRECOMP_N2[106] =  18'sd    811;
assign PRECOMP_N2[107] =  18'sd   2471;
assign PRECOMP_N2[108] =  18'sd   2433;
assign PRECOMP_N2[109] =  18'sd   1014;
assign PRECOMP_N2[110] = -18'sd    752;
assign PRECOMP_N2[111] = -18'sd   1801;
assign PRECOMP_N2[112] = -18'sd   1647;
assign PRECOMP_N2[113] = -18'sd    564;
assign PRECOMP_N2[114] =  18'sd    680;
assign PRECOMP_N2[115] =  18'sd   1340;
assign PRECOMP_N2[116] =  18'sd   1120;
assign PRECOMP_N2[117] =  18'sd    279;
assign PRECOMP_N2[118] = -18'sd    599;
assign PRECOMP_N2[119] = -18'sd    993;
assign PRECOMP_N2[120] = -18'sd    744;
assign PRECOMP_N2[121] = -18'sd     94;
assign PRECOMP_N2[122] =  18'sd    513;
assign PRECOMP_N2[123] =  18'sd    722;
assign PRECOMP_N2[124] =  18'sd    469;
assign PRECOMP_N2[125] = -18'sd     24;
assign PRECOMP_N2[126] = -18'sd    424;
assign PRECOMP_N2[127] = -18'sd    504;
assign PRECOMP_N2[128] = -18'sd    266;
assign PRECOMP_N2[129] =  18'sd     95;
assign PRECOMP_N2[130] =  18'sd    338;
assign PRECOMP_N2[131] =  18'sd    331;
assign PRECOMP_N2[132] =  18'sd    120;
assign PRECOMP_N2[133] = -18'sd    131;
assign PRECOMP_N2[134] = -18'sd    256;
assign PRECOMP_N2[135] = -18'sd    195;
assign PRECOMP_N2[136] = -18'sd     18;
assign PRECOMP_N2[137] =  18'sd    142;
assign PRECOMP_N2[138] =  18'sd    181;
assign PRECOMP_N2[139] =  18'sd     91;
assign PRECOMP_N2[140] = -18'sd     48;
assign PRECOMP_N2[141] = -18'sd    135;
assign PRECOMP_N2[142] = -18'sd    115;
assign PRECOMP_N2[143] = -18'sd     15;
assign PRECOMP_N2[144] =  18'sd     86;
assign PRECOMP_N2[145] =  18'sd    117;
assign PRECOMP_N2[146] =  18'sd     60;
assign PRECOMP_N2[147] = -18'sd     37;
assign PRECOMP_N2[148] = -18'sd    102;
assign PRECOMP_N2[149] = -18'sd     92;
assign PRECOMP_N2[150] = -18'sd     16;
assign PRECOMP_N2[151] =  18'sd     68;
assign PRECOMP_N2[152] =  18'sd    103;
assign PRECOMP_N2[153] =  18'sd     65;
assign PRECOMP_N2[154] = -18'sd     16;
assign PRECOMP_N2[155] = -18'sd     84;
assign PRECOMP_N2[156] = -18'sd     92;
assign PRECOMP_N2[157] = -18'sd     38;
assign PRECOMP_N2[158] =  18'sd     38;
assign PRECOMP_N2[159] =  18'sd     86;
assign PRECOMP_N2[160] =  18'sd     74;
assign PRECOMP_N2[161] =  18'sd     15;
assign PRECOMP_N2[162] = -18'sd     51;
assign PRECOMP_N2[163] = -18'sd     79;
assign PRECOMP_N2[164] = -18'sd     54;
assign PRECOMP_N2[165] =  18'sd      4;
assign PRECOMP_N2[166] =  18'sd     55;
assign PRECOMP_N2[167] =  18'sd     66;
assign PRECOMP_N2[168] =  18'sd     33;
assign PRECOMP_N2[169] = -18'sd     18;
assign PRECOMP_N2[170] = -18'sd     53;
assign PRECOMP_N2[171] = -18'sd     50;
assign PRECOMP_N2[172] = -18'sd     14;
assign PRECOMP_N2[173] =  18'sd     27;
assign PRECOMP_N2[174] =  18'sd     47;
assign PRECOMP_N2[175] =  18'sd     33;
assign PRECOMP_N2[176] = -18'sd      2;
assign PRECOMP_N2[177] = -18'sd     31;
assign PRECOMP_N2[178] = -18'sd     37;
assign PRECOMP_N2[179] = -18'sd     17;
assign PRECOMP_N2[180] =  18'sd     13;
assign PRECOMP_N2[181] =  18'sd     32;
assign PRECOMP_N2[182] =  18'sd     26;
assign PRECOMP_N2[183] =  18'sd      3;
assign PRECOMP_N2[184] = -18'sd     21;
assign PRECOMP_N2[185] = -18'sd     28;
assign PRECOMP_N2[186] = -18'sd     15;
assign PRECOMP_N2[187] =  18'sd      8;
assign PRECOMP_N2[188] =  18'sd     24;

