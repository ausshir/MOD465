
//RX Filter 18'sd Multiplier Coefficients (headroom)
assign coef[  0] = -18'sd    148;
assign coef[  1] = -18'sd    152;
assign coef[  2] = -18'sd     37;
assign coef[  3] =  18'sd    118;
assign coef[  4] =  18'sd    197;
assign coef[  5] =  18'sd    133;
assign coef[  6] = -18'sd     41;
assign coef[  7] = -18'sd    202;
assign coef[  8] = -18'sd    229;
assign coef[  9] = -18'sd     87;
assign coef[ 10] =  18'sd    133;
assign coef[ 11] =  18'sd    277;
assign coef[ 12] =  18'sd    232;
assign coef[ 13] =  18'sd     15;
assign coef[ 14] = -18'sd    231;
assign coef[ 15] = -18'sd    329;
assign coef[ 16] = -18'sd    199;
assign coef[ 17] =  18'sd     82;
assign coef[ 18] =  18'sd    319;
assign coef[ 19] =  18'sd    341;
assign coef[ 20] =  18'sd    120;
assign coef[ 21] = -18'sd    194;
assign coef[ 22] = -18'sd    379;
assign coef[ 23] = -18'sd    294;
assign coef[ 24] =  18'sd      7;
assign coef[ 25] =  18'sd    310;
assign coef[ 26] =  18'sd    388;
assign coef[ 27] =  18'sd    172;
assign coef[ 28] = -18'sd    185;
assign coef[ 29] = -18'sd    414;
assign coef[ 30] = -18'sd    322;
assign coef[ 31] =  18'sd     43;
assign coef[ 32] =  18'sd    413;
assign coef[ 33] =  18'sd    483;
assign coef[ 34] =  18'sd    152;
assign coef[ 35] = -18'sd    369;
assign coef[ 36] = -18'sd    684;
assign coef[ 37] = -18'sd    491;
assign coef[ 38] =  18'sd    154;
assign coef[ 39] =  18'sd    824;
assign coef[ 40] =  18'sd    988;
assign coef[ 41] =  18'sd    404;
assign coef[ 42] = -18'sd    635;
assign coef[ 43] = -18'sd   1428;
assign coef[ 44] = -18'sd   1313;
assign coef[ 45] = -18'sd    181;
assign coef[ 46] =  18'sd   1342;
assign coef[ 47] =  18'sd   2209;
assign coef[ 48] =  18'sd   1644;
assign coef[ 49] = -18'sd    239;
assign coef[ 50] = -18'sd   2350;
assign coef[ 51] = -18'sd   3217;
assign coef[ 52] = -18'sd   1964;
assign coef[ 53] =  18'sd    950;
assign coef[ 54] =  18'sd   3797;
assign coef[ 55] =  18'sd   4553;
assign coef[ 56] =  18'sd   2254;
assign coef[ 57] = -18'sd   2127;
assign coef[ 58] = -18'sd   5967;
assign coef[ 59] = -18'sd   6459;
assign coef[ 60] = -18'sd   2500;
assign coef[ 61] =  18'sd   4191;
assign coef[ 62] =  18'sd   9614;
assign coef[ 63] =  18'sd   9631;
assign coef[ 64] =  18'sd   2687;
assign coef[ 65] = -18'sd   8506;
assign coef[ 66] = -18'sd  17524;
assign coef[ 67] = -18'sd  17063;
assign coef[ 68] = -18'sd   2804;
assign coef[ 69] =  18'sd  23719;
assign coef[ 70] =  18'sd  54919;
assign coef[ 71] =  18'sd  79992;
assign coef[ 72] =  18'sd  89579;
