
//TX Filter 18'sd Multiplier Coefficients (headroom)
assign coef[  0] = -18'sd     50;
assign coef[  1] = -18'sd     87;
assign coef[  2] = -18'sd     60;
assign coef[  3] =  18'sd     18;
assign coef[  4] =  18'sd     96;
assign coef[  5] =  18'sd    111;
assign coef[  6] =  18'sd     40;
assign coef[  7] = -18'sd     79;
assign coef[  8] = -18'sd    160;
assign coef[  9] = -18'sd    131;
assign coef[ 10] =  18'sd      8;
assign coef[ 11] =  18'sd    172;
assign coef[ 12] =  18'sd    241;
assign coef[ 13] =  18'sd    139;
assign coef[ 14] = -18'sd     93;
assign coef[ 15] = -18'sd    308;
assign coef[ 16] = -18'sd    340;
assign coef[ 17] = -18'sd    127;
assign coef[ 18] =  18'sd    228;
assign coef[ 19] =  18'sd    493;
assign coef[ 20] =  18'sd    456;
assign coef[ 21] =  18'sd     82;
assign coef[ 22] = -18'sd    428;
assign coef[ 23] = -18'sd    737;
assign coef[ 24] = -18'sd    586;
assign coef[ 25] =  18'sd      9;
assign coef[ 26] =  18'sd    712;
assign coef[ 27] =  18'sd   1053;
assign coef[ 28] =  18'sd    726;
assign coef[ 29] = -18'sd    165;
assign coef[ 30] = -18'sd   1104;
assign coef[ 31] = -18'sd   1454;
assign coef[ 32] = -18'sd    870;
assign coef[ 33] =  18'sd    411;
assign coef[ 34] =  18'sd   1638;
assign coef[ 35] =  18'sd   1964;
assign coef[ 36] =  18'sd   1014;
assign coef[ 37] = -18'sd    788;
assign coef[ 38] = -18'sd   2369;
assign coef[ 39] = -18'sd   2623;
assign coef[ 40] = -18'sd   1150;
assign coef[ 41] =  18'sd   1360;
assign coef[ 42] =  18'sd   3400;
assign coef[ 43] =  18'sd   3514;
assign coef[ 44] =  18'sd   1273;
assign coef[ 45] = -18'sd   2257;
assign coef[ 46] = -18'sd   4948;
assign coef[ 47] = -18'sd   4822;
assign coef[ 48] = -18'sd   1375;
assign coef[ 49] =  18'sd   3793;
assign coef[ 50] =  18'sd   7585;
assign coef[ 51] =  18'sd   7081;
assign coef[ 52] =  18'sd   1453;
assign coef[ 53] = -18'sd   6996;
assign coef[ 54] = -18'sd  13415;
assign coef[ 55] = -18'sd  12554;
assign coef[ 56] = -18'sd   1501;
assign coef[ 57] =  18'sd  18381;
assign coef[ 58] =  18'sd  41444;
assign coef[ 59] =  18'sd  59844;
assign coef[ 60] =  18'sd  66857;
